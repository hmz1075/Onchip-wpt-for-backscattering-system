magic
tech sky130A
timestamp 1634733432
<< metal5 >>
rect 394000 1624000 683000 1631000
rect 394000 1449000 401000 1624000
rect 405000 1613000 672000 1620000
rect 405000 1460000 412000 1613000
rect 419500 1602000 661000 1609000
rect 654000 1460000 661000 1602000
rect 405000 1453000 661000 1460000
rect 665000 1449000 672000 1613000
rect 394000 1442000 672000 1449000
rect 676000 1438000 683000 1624000
rect 397000 1431000 683000 1438000
<< end >>
