magic
tech sky130A
magscale 1 2
timestamp 1634285219
<< error_p >>
rect -31 8081 31 8087
rect -31 8047 -19 8081
rect -31 8041 31 8047
rect -31 -8047 31 -8041
rect -31 -8081 -19 -8047
rect -31 -8087 31 -8081
<< nwell >>
rect -231 -8219 231 8219
<< pmos >>
rect -35 -8000 35 8000
<< pdiff >>
rect -93 7988 -35 8000
rect -93 -7988 -81 7988
rect -47 -7988 -35 7988
rect -93 -8000 -35 -7988
rect 35 7988 93 8000
rect 35 -7988 47 7988
rect 81 -7988 93 7988
rect 35 -8000 93 -7988
<< pdiffc >>
rect -81 -7988 -47 7988
rect 47 -7988 81 7988
<< nsubdiff >>
rect -195 8149 -99 8183
rect 99 8149 195 8183
rect -195 8087 -161 8149
rect 161 8087 195 8149
rect -195 -8149 -161 -8087
rect 161 -8149 195 -8087
rect -195 -8183 -99 -8149
rect 99 -8183 195 -8149
<< nsubdiffcont >>
rect -99 8149 99 8183
rect -195 -8087 -161 8087
rect 161 -8087 195 8087
rect -99 -8183 99 -8149
<< poly >>
rect -35 8081 35 8097
rect -35 8047 -19 8081
rect 19 8047 35 8081
rect -35 8000 35 8047
rect -35 -8047 35 -8000
rect -35 -8081 -19 -8047
rect 19 -8081 35 -8047
rect -35 -8097 35 -8081
<< polycont >>
rect -19 8047 19 8081
rect -19 -8081 19 -8047
<< locali >>
rect -195 8149 -99 8183
rect 99 8149 195 8183
rect -195 8087 -161 8149
rect 161 8087 195 8149
rect -35 8047 -19 8081
rect 19 8047 35 8081
rect -81 7988 -47 8004
rect -81 -8004 -47 -7988
rect 47 7988 81 8004
rect 47 -8004 81 -7988
rect -35 -8081 -19 -8047
rect 19 -8081 35 -8047
rect -195 -8149 -161 -8087
rect 161 -8149 195 -8087
rect -195 -8183 -99 -8149
rect 99 -8183 195 -8149
<< viali >>
rect -19 8047 19 8081
rect -81 -7988 -47 7988
rect 47 -7988 81 7988
rect -19 -8081 19 -8047
<< metal1 >>
rect -31 8081 31 8087
rect -31 8047 -19 8081
rect 19 8047 31 8081
rect -31 8041 31 8047
rect -87 7988 -41 8000
rect -87 -7988 -81 7988
rect -47 -7988 -41 7988
rect -87 -8000 -41 -7988
rect 41 7988 87 8000
rect 41 -7988 47 7988
rect 81 -7988 87 7988
rect 41 -8000 87 -7988
rect -31 -8047 31 -8041
rect -31 -8081 -19 -8047
rect 19 -8081 31 -8047
rect -31 -8087 31 -8081
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -178 -8166 178 8166
string parameters w 80 l 0.35 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
