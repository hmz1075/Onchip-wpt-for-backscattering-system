magic
tech sky130A
magscale 1 2
timestamp 1634293569
<< nwell >>
rect 3788 2096 3822 2876
rect 14120 2390 14154 2930
rect 3872 2262 3922 2312
<< pwell >>
rect 9086 1926 9840 2018
rect 4852 1788 4912 1860
rect 8968 1786 9028 1858
rect 9880 1778 9952 1862
rect 4772 1516 4806 1684
rect 5160 1418 6130 1772
rect 9086 1504 9120 1672
rect 9806 1496 9840 1664
rect 14120 1484 14154 1652
rect 4854 1334 4914 1406
rect 8970 1334 9030 1406
<< psubdiff >>
rect 4772 1516 4806 1684
rect 9086 1504 9120 1672
rect 9806 1496 9840 1664
rect 14120 1484 14154 1652
<< nsubdiff >>
rect 3788 2096 3822 2876
rect 14120 2390 14154 2930
<< poly >>
rect 3872 2262 3922 2312
rect 4852 1788 4912 1860
rect 8968 1786 9028 1858
rect 9880 1778 9952 1862
rect 4854 1334 4914 1406
rect 8970 1334 9030 1406
<< locali >>
rect 3788 2136 3822 2876
rect 4034 2794 4282 2938
rect 4088 2334 4336 2478
rect 14120 2390 14154 2930
rect 3788 2096 3796 2136
rect 9086 1926 9840 2018
rect 4772 1516 4806 1684
rect 9086 1504 9120 1672
rect 9806 1496 9840 1664
rect 11718 1636 12618 1772
rect 14120 1484 14154 1652
rect 5416 736 6316 872
<< viali >>
rect 3796 2096 3858 2136
rect 9180 2080 9744 2120
rect 3794 618 3864 652
rect 8978 632 9024 694
<< metal1 >>
rect 3850 2776 3934 2794
rect 3850 2710 3864 2776
rect 3932 2710 3934 2776
rect 14008 2714 14062 2778
rect 3850 2692 3934 2710
rect 5100 2684 5812 2688
rect 5100 2632 5108 2684
rect 5800 2632 5812 2684
rect 5100 2608 5812 2632
rect 3862 2314 3932 2328
rect 3862 2262 3872 2314
rect 3928 2262 3932 2314
rect 3862 2252 3932 2262
rect 14010 2254 14064 2318
rect 7234 2228 7946 2230
rect 3792 2158 3886 2178
rect 3790 2136 3886 2158
rect 3790 2096 3796 2136
rect 3858 2096 3886 2136
rect 7234 2172 7252 2228
rect 7926 2172 7946 2228
rect 7234 2128 7946 2172
rect 3790 1862 3886 2096
rect 9164 2120 9760 2126
rect 9164 2080 9180 2120
rect 9744 2080 9760 2120
rect 5094 1936 5816 1950
rect 5094 1876 5100 1936
rect 5810 1876 5816 1936
rect 5094 1872 5102 1876
rect 5808 1872 5816 1876
rect 5094 1870 5816 1872
rect 9164 1862 9760 2080
rect 3790 1860 4908 1862
rect 3790 1788 4912 1860
rect 3790 1786 4908 1788
rect 3790 964 3886 1786
rect 8974 1784 9950 1862
rect 10614 1826 10630 1882
rect 11404 1826 11426 1882
rect 10614 1820 11426 1826
rect 14010 1794 14064 1858
rect 9164 1782 9760 1784
rect 6080 1772 6130 1774
rect 5182 1764 6130 1772
rect 5182 1682 5198 1764
rect 6108 1682 6130 1764
rect 5182 1678 5200 1682
rect 6092 1678 6130 1682
rect 5182 1654 6130 1678
rect 5182 1648 6102 1654
rect 5152 1512 6136 1522
rect 5152 1424 5164 1512
rect 6120 1424 6136 1512
rect 10602 1488 11454 1502
rect 4854 1334 4914 1406
rect 6338 1382 6366 1438
rect 6916 1382 6928 1438
rect 10602 1432 10616 1488
rect 11428 1432 11454 1488
rect 6338 1372 6928 1382
rect 8974 1402 9950 1404
rect 7222 1362 7978 1378
rect 4028 1308 4294 1330
rect 4028 1222 4044 1308
rect 4256 1304 4294 1308
rect 4256 1222 5162 1304
rect 7222 1298 7238 1362
rect 7966 1298 7978 1362
rect 8974 1334 9214 1402
rect 9694 1334 9950 1402
rect 14010 1332 14064 1396
rect 7222 1296 7978 1298
rect 11690 1238 11712 1282
rect 12594 1238 12610 1282
rect 11690 1226 12610 1238
rect 4028 1212 5162 1222
rect 4028 1210 4294 1212
rect 6340 1044 6914 1064
rect 6340 994 6354 1044
rect 6900 994 6914 1044
rect 3790 880 4914 964
rect 3790 658 3886 880
rect 8978 704 9034 960
rect 8960 694 9054 704
rect 3786 652 3894 658
rect 3786 618 3794 652
rect 3864 618 3894 652
rect 3786 586 3894 618
rect 8960 632 8978 694
rect 9024 632 9054 694
rect 8960 608 9054 632
rect 11674 580 12618 592
rect 11674 524 11696 580
rect 12580 524 12618 580
rect 11674 522 12618 524
rect 3874 490 3944 494
rect 3874 434 3882 490
rect 3936 434 3944 490
rect 3874 430 3944 434
rect 9206 460 9698 472
rect 9206 392 9214 460
rect 9694 392 9698 460
rect 14012 428 14066 492
<< via1 >>
rect 3864 2710 3932 2776
rect 5108 2632 5800 2684
rect 3872 2262 3928 2314
rect 7252 2172 7926 2228
rect 5100 1876 5810 1936
rect 5102 1872 5808 1876
rect 10630 1826 11404 1888
rect 5198 1682 6108 1764
rect 5200 1678 6092 1682
rect 5164 1418 6120 1512
rect 6366 1382 6916 1438
rect 10616 1428 11428 1488
rect 4044 1222 4256 1308
rect 7238 1298 7966 1362
rect 9214 1334 9694 1402
rect 11712 1238 12594 1304
rect 6354 986 6900 1044
rect 11696 524 12580 580
rect 3882 434 3936 490
rect 9214 392 9694 460
<< metal2 >>
rect 3846 2780 3940 2794
rect 3846 2710 3864 2780
rect 3934 2714 3940 2780
rect 3932 2710 3940 2714
rect 3846 2686 3940 2710
rect 5092 2684 5824 2698
rect 5092 2632 5108 2684
rect 5800 2632 5824 2684
rect 5092 2344 5824 2632
rect 3866 2314 5824 2344
rect 3866 2262 3872 2314
rect 3928 2262 5824 2314
rect 3866 2226 5824 2262
rect 3954 2220 5824 2226
rect 5092 1936 5824 2220
rect 5092 1876 5100 1936
rect 5810 1876 5824 1936
rect 5092 1872 5102 1876
rect 5808 1872 5824 1876
rect 5092 1870 5824 1872
rect 7214 2228 7992 2234
rect 7214 2172 7252 2228
rect 7926 2172 7992 2228
rect 5160 1764 6130 1772
rect 5160 1682 5198 1764
rect 6108 1682 6130 1764
rect 5160 1678 5200 1682
rect 6092 1678 6130 1682
rect 5160 1542 6130 1678
rect 5164 1512 6130 1542
rect 6120 1418 6130 1512
rect 6338 1438 6932 1444
rect 5164 1394 5326 1418
rect 6338 1382 6366 1438
rect 6916 1382 6932 1438
rect 3954 1326 4292 1330
rect 3866 1316 4292 1326
rect 3866 1226 3886 1316
rect 3942 1308 4292 1316
rect 3942 1226 4044 1308
rect 3866 1222 4044 1226
rect 4256 1222 4292 1308
rect 3866 1210 4292 1222
rect 3870 494 3936 1210
rect 6338 1044 6932 1382
rect 7214 1362 7992 2172
rect 10606 1888 11466 1896
rect 10606 1826 10630 1888
rect 11404 1826 11466 1888
rect 10606 1488 11466 1826
rect 10606 1428 10616 1488
rect 11428 1428 11466 1488
rect 10606 1420 11466 1428
rect 7214 1298 7238 1362
rect 7966 1298 7992 1362
rect 7214 1290 7992 1298
rect 9206 1402 9706 1404
rect 9206 1334 9214 1402
rect 9694 1334 9706 1402
rect 6338 986 6354 1044
rect 6900 986 6932 1044
rect 6338 980 6932 986
rect 9206 598 9706 1334
rect 3870 490 3944 494
rect 3870 434 3882 490
rect 3936 434 3944 490
rect 3870 430 3944 434
rect 9204 460 9706 598
rect 11684 1304 12628 1312
rect 11684 1238 11712 1304
rect 12594 1238 12628 1304
rect 11684 580 12628 1238
rect 11684 524 11696 580
rect 12580 524 12628 580
rect 11684 514 12628 524
rect 9204 392 9214 460
rect 9694 392 9706 460
rect 9204 386 9706 392
rect 9204 -276 9704 386
<< via2 >>
rect 3864 2776 3934 2780
rect 3864 2714 3932 2776
rect 3932 2714 3934 2776
rect 3886 1226 3942 1316
<< metal3 >>
rect 3836 2780 3950 2804
rect 3836 2714 3864 2780
rect 3934 2714 3950 2780
rect 3836 2668 3950 2714
rect 3878 1316 3948 2668
rect 3878 1226 3886 1316
rect 3942 1226 3948 1316
rect 3878 1208 3948 1226
use sky130_fd_pr__nfet_01v8_lvt_8K7EBA  sky130_fd_pr__nfet_01v8_lvt_8K7EBA_1
timestamp 1634293406
transform 0 1 6946 -1 0 925
box -231 -2210 231 2210
use sky130_fd_pr__nfet_01v8_lvt_8K7EBA  sky130_fd_pr__nfet_01v8_lvt_8K7EBA_0
timestamp 1634293406
transform 0 -1 6946 -1 0 1369
box -231 -2210 231 2210
use sky130_fd_pr__nfet_01v8_lvt_8K7EBA  sky130_fd_pr__nfet_01v8_lvt_8K7EBA_3
timestamp 1634293406
transform 0 1 6946 -1 0 1823
box -231 -2210 231 2210
use sky130_fd_pr__nfet_01v8_lvt_8K7EBA  sky130_fd_pr__nfet_01v8_lvt_8K7EBA_2
timestamp 1634293406
transform 0 1 11980 -1 0 1367
box -231 -2210 231 2210
use sky130_fd_pr__nfet_01v8_lvt_8K7EBA  sky130_fd_pr__nfet_01v8_lvt_8K7EBA_4
timestamp 1634293406
transform 0 1 11980 -1 0 1825
box -231 -2210 231 2210
use sky130_fd_pr__pfet_01v8_lvt_4QC8GG  sky130_fd_pr__pfet_01v8_lvt_4QC8GG_0
timestamp 1634206901
transform 0 1 8971 -1 0 2287
box -231 -5219 231 5219
use sky130_fd_pr__pfet_01v8_lvt_4QC8GG  sky130_fd_pr__pfet_01v8_lvt_4QC8GG_1
timestamp 1634206901
transform 0 1 8971 -1 0 2745
box -231 -5219 231 5219
use sky130_fd_pr__pfet_01v8_lvt_4QC8GG  sky130_fd_pr__pfet_01v8_lvt_4QC8GG_2
timestamp 1634206901
transform 0 1 8973 -1 0 459
box -231 -5219 231 5219
<< labels >>
rlabel metal1 3816 1492 3816 1492 1 VIN-
rlabel metal2 12062 882 12062 882 1 VOUT
rlabel locali 14138 1550 14138 1550 1 VSS
rlabel metal2 9454 -218 9454 -218 1 VINp
<< end >>
