magic
tech sky130A
magscale 1 2
timestamp 1634295700
<< locali >>
rect -18 16312 9156 16348
rect -18 -18 9150 18
<< metal1 >>
rect 144 16252 9216 16344
rect 142 16240 9216 16252
rect 142 16214 8992 16240
rect 142 16208 672 16214
rect -238 16168 132 16172
rect 946 16168 1050 16176
rect -238 16116 34 16168
rect 94 16116 132 16168
rect -238 16100 132 16116
rect 482 16164 586 16168
rect 482 16112 490 16164
rect 550 16112 586 16164
rect 946 16116 952 16168
rect 1012 16116 1050 16168
rect 946 16112 1050 16116
rect 1402 16164 1506 16172
rect 1402 16112 1410 16164
rect 1470 16112 1506 16164
rect 1868 16170 1972 16176
rect 1868 16118 1874 16170
rect 1934 16118 1972 16170
rect 1868 16112 1972 16118
rect 2328 16174 2432 16180
rect 2328 16122 2332 16174
rect 2392 16122 2432 16174
rect 2328 16116 2432 16122
rect 2796 16174 2900 16182
rect 2796 16122 2802 16174
rect 2862 16122 2900 16174
rect 3254 16176 3358 16186
rect 3254 16124 3260 16176
rect 3320 16124 3358 16176
rect 3254 16122 3358 16124
rect 3716 16176 3820 16184
rect 3716 16124 3724 16176
rect 3784 16124 3820 16176
rect 2796 16118 2900 16122
rect 3716 16120 3820 16124
rect 4178 16176 4282 16184
rect 4178 16124 4186 16176
rect 4246 16124 4282 16176
rect 4178 16120 4282 16124
rect 4640 16176 4744 16182
rect 4640 16124 4648 16176
rect 4708 16124 4744 16176
rect 4640 16118 4744 16124
rect 5100 16176 5204 16186
rect 5100 16124 5108 16176
rect 5168 16124 5204 16176
rect 5100 16122 5204 16124
rect 5564 16176 5668 16184
rect 5564 16124 5572 16176
rect 5632 16124 5668 16176
rect 5564 16120 5668 16124
rect 6026 16180 6130 16186
rect 6026 16128 6032 16180
rect 6092 16128 6130 16180
rect 6026 16122 6130 16128
rect 6484 16174 6588 16184
rect 6484 16122 6498 16174
rect 6558 16122 6588 16174
rect 6948 16176 7052 16186
rect 6948 16124 6956 16176
rect 7016 16124 7052 16176
rect 6948 16122 7052 16124
rect 7408 16178 7512 16186
rect 7408 16126 7422 16178
rect 7482 16126 7512 16178
rect 7408 16122 7512 16126
rect 7872 16178 7976 16186
rect 7872 16126 7884 16178
rect 7944 16126 7976 16178
rect 7872 16122 7976 16126
rect 8334 16178 8438 16186
rect 8334 16126 8344 16178
rect 8404 16126 8438 16178
rect 8334 16122 8438 16126
rect 8794 16172 8898 16180
rect 6484 16120 6588 16122
rect 8794 16120 8806 16172
rect 8866 16120 8898 16172
rect 8794 16116 8898 16120
rect 482 16104 586 16112
rect 1402 16108 1506 16112
rect 224 230 340 236
rect 224 176 272 230
rect 328 176 340 230
rect 224 162 340 176
rect 684 232 800 240
rect 684 178 730 232
rect 786 178 800 232
rect 684 166 800 178
rect 1142 236 1258 240
rect 1142 182 1196 236
rect 1252 182 1258 236
rect 1142 166 1258 182
rect 1606 234 1722 240
rect 1606 180 1652 234
rect 1708 180 1722 234
rect 1606 166 1722 180
rect 2066 232 2182 240
rect 2066 178 2112 232
rect 2168 178 2182 232
rect 2066 166 2182 178
rect 2528 236 2644 240
rect 2528 182 2580 236
rect 2636 182 2644 236
rect 2528 166 2644 182
rect 2990 230 3106 240
rect 2990 176 3044 230
rect 3100 176 3106 230
rect 2990 166 3106 176
rect 3452 232 3568 240
rect 3452 178 3506 232
rect 3562 178 3568 232
rect 3452 166 3568 178
rect 3914 234 4030 240
rect 3914 180 3966 234
rect 4022 180 4030 234
rect 3914 166 4030 180
rect 4376 234 4492 240
rect 4376 180 4426 234
rect 4482 180 4492 234
rect 4376 166 4492 180
rect 4840 230 4956 240
rect 4840 176 4886 230
rect 4942 176 4956 230
rect 4840 166 4956 176
rect 5302 232 5418 240
rect 5302 178 5350 232
rect 5406 178 5418 232
rect 5302 166 5418 178
rect 5762 230 5878 236
rect 5762 176 5812 230
rect 5868 176 5878 230
rect 5762 162 5878 176
rect 6224 232 6340 240
rect 6224 178 6274 232
rect 6330 178 6340 232
rect 6224 166 6340 178
rect 6688 234 6804 242
rect 6688 180 6740 234
rect 6796 180 6804 234
rect 6688 168 6804 180
rect 7150 234 7266 238
rect 7150 180 7200 234
rect 7256 180 7266 234
rect 7150 164 7266 180
rect 7612 234 7728 238
rect 7612 180 7662 234
rect 7718 180 7728 234
rect 7612 164 7728 180
rect 8070 232 8186 238
rect 8070 178 8124 232
rect 8180 178 8186 232
rect 8070 164 8186 178
rect 8536 232 8652 240
rect 8536 178 8584 232
rect 8640 178 8652 232
rect 8536 166 8652 178
rect 8996 232 9112 238
rect 8996 178 9054 232
rect 9110 178 9112 232
rect 8996 164 9112 178
rect 140 -278 9006 126
<< via1 >>
rect 34 16116 94 16168
rect 490 16112 550 16164
rect 952 16116 1012 16168
rect 1410 16112 1470 16164
rect 1874 16118 1934 16170
rect 2332 16122 2392 16174
rect 2802 16122 2862 16174
rect 3260 16124 3320 16176
rect 3724 16124 3784 16176
rect 4186 16124 4246 16176
rect 4648 16124 4708 16176
rect 5108 16124 5168 16176
rect 5572 16124 5632 16176
rect 6032 16128 6092 16180
rect 6498 16122 6558 16174
rect 6956 16124 7016 16176
rect 7422 16126 7482 16178
rect 7884 16126 7944 16178
rect 8344 16126 8404 16178
rect 8806 16120 8866 16172
rect 272 176 328 230
rect 730 178 786 232
rect 1196 182 1252 236
rect 1652 180 1708 234
rect 2112 178 2168 232
rect 2580 182 2636 236
rect 3044 176 3100 230
rect 3506 178 3562 232
rect 3966 180 4022 234
rect 4426 180 4482 234
rect 4886 176 4942 230
rect 5350 178 5406 232
rect 5812 176 5868 230
rect 6274 178 6330 232
rect 6740 180 6796 234
rect 7200 180 7256 234
rect 7662 180 7718 234
rect 8124 178 8180 232
rect 8584 178 8640 232
rect 9054 178 9110 232
<< metal2 >>
rect 22 16176 6032 16180
rect 22 16174 3260 16176
rect 22 16170 2332 16174
rect 22 16168 1874 16170
rect 22 16116 34 16168
rect 94 16164 952 16168
rect 94 16116 490 16164
rect 22 16112 490 16116
rect 550 16116 952 16164
rect 1012 16164 1874 16168
rect 1012 16116 1410 16164
rect 550 16112 1410 16116
rect 1470 16118 1874 16164
rect 1934 16122 2332 16170
rect 2392 16122 2802 16174
rect 2862 16124 3260 16174
rect 3320 16124 3724 16176
rect 3784 16124 4186 16176
rect 4246 16124 4648 16176
rect 4708 16124 5108 16176
rect 5168 16124 5572 16176
rect 5632 16128 6032 16176
rect 6092 16178 8918 16180
rect 6092 16176 7422 16178
rect 6092 16174 6956 16176
rect 6092 16128 6498 16174
rect 5632 16124 6498 16128
rect 2862 16122 6498 16124
rect 6558 16124 6956 16174
rect 7016 16126 7422 16176
rect 7482 16126 7884 16178
rect 7944 16126 8344 16178
rect 8404 16172 8918 16178
rect 8404 16126 8806 16172
rect 7016 16124 8806 16126
rect 6558 16122 8806 16124
rect 1934 16120 8806 16122
rect 8866 16120 8918 16172
rect 1934 16118 8918 16120
rect 1470 16112 8918 16118
rect 22 16102 8918 16112
rect -154 236 9114 240
rect -154 232 1196 236
rect -154 230 730 232
rect -154 176 272 230
rect 328 178 730 230
rect 786 182 1196 232
rect 1252 234 2580 236
rect 1252 182 1652 234
rect 786 180 1652 182
rect 1708 232 2580 234
rect 1708 180 2112 232
rect 786 178 2112 180
rect 2168 182 2580 232
rect 2636 234 9114 236
rect 2636 232 3966 234
rect 2636 230 3506 232
rect 2636 182 3044 230
rect 2168 178 3044 182
rect 328 176 3044 178
rect 3100 178 3506 230
rect 3562 180 3966 232
rect 4022 180 4426 234
rect 4482 232 6740 234
rect 4482 230 5350 232
rect 4482 180 4886 230
rect 3562 178 4886 180
rect 3100 176 4886 178
rect 4942 178 5350 230
rect 5406 230 6274 232
rect 5406 178 5812 230
rect 4942 176 5812 178
rect 5868 178 6274 230
rect 6330 180 6740 232
rect 6796 180 7200 234
rect 7256 180 7662 234
rect 7718 232 9114 234
rect 7718 180 8124 232
rect 6330 178 8124 180
rect 8180 178 8584 232
rect 8640 178 9054 232
rect 9110 178 9114 232
rect 5868 176 9114 178
rect -154 166 9114 176
rect -154 162 342 166
use sky130_fd_pr__pfet_01v8_lvt_4QDPGG  sky130_fd_pr__pfet_01v8_lvt_4QDPGG_0
array 19 0 462 0 0 16438
timestamp 1634285219
transform 1 0 178 0 1 8166
box -231 -8219 231 8219
<< labels >>
rlabel metal1 -216 16116 -216 16116 1 D
rlabel metal2 -132 200 -132 200 1 S
rlabel locali 9120 -6 9120 -6 1 B
rlabel metal1 504 -162 504 -162 1 G
<< end >>
