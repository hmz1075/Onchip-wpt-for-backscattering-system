magic
tech sky130A
magscale 1 2
timestamp 1634725508
<< metal1 >>
rect -480 38320 948 38438
rect -480 37928 -288 38320
rect 546 37928 948 38320
rect -480 37872 948 37928
rect -480 37868 -396 37872
rect 848 37792 948 37872
rect 882 37746 948 37792
rect 882 37730 904 37746
rect 936 37556 948 37746
rect 17684 520 18170 594
rect 17684 514 18210 520
rect 17435 446 18210 514
rect 17435 156 17834 446
rect 18096 156 18210 446
rect 17435 56 18210 156
rect 17714 42 18210 56
<< via1 >>
rect -288 37928 546 38320
rect 17834 156 18096 446
<< metal2 >>
rect -390 39902 590 40110
rect -390 39186 -278 39902
rect 462 39186 590 39902
rect -390 38592 590 39186
rect -396 38320 660 38592
rect -396 37928 -288 38320
rect 546 37928 660 38320
rect -396 37894 660 37928
rect -390 37890 -246 37894
rect 480 37890 590 37894
rect 17714 446 18210 520
rect 17714 156 17834 446
rect 18096 156 18210 446
rect 17714 42 18210 156
rect 17770 30 18164 42
<< via2 >>
rect -278 39186 462 39902
rect 17834 156 18096 446
<< metal3 >>
rect -390 39902 624 45240
rect -390 39186 -278 39902
rect 462 39186 624 39902
rect -390 38960 624 39186
rect 17714 446 18210 520
rect 17714 156 17834 446
rect 18096 156 18210 446
rect 17714 42 18210 156
rect 17770 30 18164 42
<< via3 >>
rect 17834 156 18096 446
<< metal4 >>
rect 17760 520 18152 41498
rect 17714 446 18210 520
rect 17714 156 17834 446
rect 18096 156 18210 446
rect 17714 42 18210 156
use cap107_layout  cap107_layout_0
timestamp 1634724870
transform 1 0 30066 0 1 87546
box -87990 -83672 8182 10526
use FINAL  FINAL_0
timestamp 1634546801
transform 1 0 2 0 1 2
box -2 -2 136810 98784
<< labels >>
rlabel metal2 -72 38660 -72 38660 1 VINN
rlabel metal4 17974 40444 17974 40444 1 VINP
<< end >>
