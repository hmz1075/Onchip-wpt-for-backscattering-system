magic
tech sky130A
magscale 1 2
timestamp 1634546801
<< error_p >>
rect -18467 18370 -18247 24190
rect -24306 18230 -18247 18370
rect -18227 18370 -18007 24190
rect -12388 18370 -12168 24190
rect -18227 18230 -12168 18370
rect -12148 18370 -11928 24190
rect -6309 18370 -6089 24190
rect -12148 18230 -6089 18370
rect -6069 18370 -5849 24190
rect -230 18370 -10 24190
rect -6069 18230 -10 18370
rect 10 18370 230 24190
rect 5849 18370 6069 24190
rect 10 18230 6069 18370
rect 6089 18370 6309 24190
rect 11928 18370 12148 24190
rect 6089 18230 12148 18370
rect 12168 18370 12388 24190
rect 18007 18370 18227 24190
rect 12168 18230 18227 18370
rect 18247 18370 18467 24190
rect 18247 18230 24306 18370
rect -24306 17990 -18247 18130
rect -18467 12310 -18247 17990
rect -24306 12170 -18247 12310
rect -18227 17990 -12168 18130
rect -18227 12310 -18007 17990
rect -12388 12310 -12168 17990
rect -18227 12170 -12168 12310
rect -12148 17990 -6089 18130
rect -12148 12310 -11928 17990
rect -6309 12310 -6089 17990
rect -12148 12170 -6089 12310
rect -6069 17990 -10 18130
rect -6069 12310 -5849 17990
rect -230 12310 -10 17990
rect -6069 12170 -10 12310
rect 10 17990 6069 18130
rect 10 12310 230 17990
rect 5849 12310 6069 17990
rect 10 12170 6069 12310
rect 6089 17990 12148 18130
rect 6089 12310 6309 17990
rect 11928 12310 12148 17990
rect 6089 12170 12148 12310
rect 12168 17990 18227 18130
rect 12168 12310 12388 17990
rect 18007 12310 18227 17990
rect 12168 12170 18227 12310
rect 18247 17990 24306 18130
rect 18247 12310 18467 17990
rect 18247 12170 24306 12310
rect -24306 11930 -18247 12070
rect -18467 6250 -18247 11930
rect -24306 6110 -18247 6250
rect -18227 11930 -12168 12070
rect -18227 6250 -18007 11930
rect -12388 6250 -12168 11930
rect -18227 6110 -12168 6250
rect -12148 11930 -6089 12070
rect -12148 6250 -11928 11930
rect -6309 6250 -6089 11930
rect -12148 6110 -6089 6250
rect -6069 11930 -10 12070
rect -6069 6250 -5849 11930
rect -230 6250 -10 11930
rect -6069 6110 -10 6250
rect 10 11930 6069 12070
rect 10 6250 230 11930
rect 5849 6250 6069 11930
rect 10 6110 6069 6250
rect 6089 11930 12148 12070
rect 6089 6250 6309 11930
rect 11928 6250 12148 11930
rect 6089 6110 12148 6250
rect 12168 11930 18227 12070
rect 12168 6250 12388 11930
rect 18007 6250 18227 11930
rect 12168 6110 18227 6250
rect 18247 11930 24306 12070
rect 18247 6250 18467 11930
rect 18247 6110 24306 6250
rect -24306 5870 -18247 6010
rect -18467 190 -18247 5870
rect -24306 50 -18247 190
rect -18227 5870 -12168 6010
rect -18227 190 -18007 5870
rect -12388 190 -12168 5870
rect -18227 50 -12168 190
rect -12148 5870 -6089 6010
rect -12148 190 -11928 5870
rect -6309 190 -6089 5870
rect -12148 50 -6089 190
rect -6069 5870 -10 6010
rect -6069 190 -5849 5870
rect -230 190 -10 5870
rect -6069 50 -10 190
rect 10 5870 6069 6010
rect 10 190 230 5870
rect 5849 190 6069 5870
rect 10 50 6069 190
rect 6089 5870 12148 6010
rect 6089 190 6309 5870
rect 11928 190 12148 5870
rect 6089 50 12148 190
rect 12168 5870 18227 6010
rect 12168 190 12388 5870
rect 18007 190 18227 5870
rect 12168 50 18227 190
rect 18247 5870 24306 6010
rect 18247 190 18467 5870
rect 18247 50 24306 190
rect -24306 -190 -18247 -50
rect -18467 -5870 -18247 -190
rect -24306 -6010 -18247 -5870
rect -18227 -190 -12168 -50
rect -18227 -5870 -18007 -190
rect -12388 -5870 -12168 -190
rect -18227 -6010 -12168 -5870
rect -12148 -190 -6089 -50
rect -12148 -5870 -11928 -190
rect -6309 -5870 -6089 -190
rect -12148 -6010 -6089 -5870
rect -6069 -190 -10 -50
rect -6069 -5870 -5849 -190
rect -230 -5870 -10 -190
rect -6069 -6010 -10 -5870
rect 10 -190 6069 -50
rect 10 -5870 230 -190
rect 5849 -5870 6069 -190
rect 10 -6010 6069 -5870
rect 6089 -190 12148 -50
rect 6089 -5870 6309 -190
rect 11928 -5870 12148 -190
rect 6089 -6010 12148 -5870
rect 12168 -190 18227 -50
rect 12168 -5870 12388 -190
rect 18007 -5870 18227 -190
rect 12168 -6010 18227 -5870
rect 18247 -190 24306 -50
rect 18247 -5870 18467 -190
rect 18247 -6010 24306 -5870
rect -24306 -6250 -18247 -6110
rect -18467 -11930 -18247 -6250
rect -24306 -12070 -18247 -11930
rect -18227 -6250 -12168 -6110
rect -18227 -11930 -18007 -6250
rect -12388 -11930 -12168 -6250
rect -18227 -12070 -12168 -11930
rect -12148 -6250 -6089 -6110
rect -12148 -11930 -11928 -6250
rect -6309 -11930 -6089 -6250
rect -12148 -12070 -6089 -11930
rect -6069 -6250 -10 -6110
rect -6069 -11930 -5849 -6250
rect -230 -11930 -10 -6250
rect -6069 -12070 -10 -11930
rect 10 -6250 6069 -6110
rect 10 -11930 230 -6250
rect 5849 -11930 6069 -6250
rect 10 -12070 6069 -11930
rect 6089 -6250 12148 -6110
rect 6089 -11930 6309 -6250
rect 11928 -11930 12148 -6250
rect 6089 -12070 12148 -11930
rect 12168 -6250 18227 -6110
rect 12168 -11930 12388 -6250
rect 18007 -11930 18227 -6250
rect 12168 -12070 18227 -11930
rect 18247 -6250 24306 -6110
rect 18247 -11930 18467 -6250
rect 18247 -12070 24306 -11930
rect -24306 -12310 -18247 -12170
rect -18467 -17990 -18247 -12310
rect -24306 -18130 -18247 -17990
rect -18227 -12310 -12168 -12170
rect -18227 -17990 -18007 -12310
rect -12388 -17990 -12168 -12310
rect -18227 -18130 -12168 -17990
rect -12148 -12310 -6089 -12170
rect -12148 -17990 -11928 -12310
rect -6309 -17990 -6089 -12310
rect -12148 -18130 -6089 -17990
rect -6069 -12310 -10 -12170
rect -6069 -17990 -5849 -12310
rect -230 -17990 -10 -12310
rect -6069 -18130 -10 -17990
rect 10 -12310 6069 -12170
rect 10 -17990 230 -12310
rect 5849 -17990 6069 -12310
rect 10 -18130 6069 -17990
rect 6089 -12310 12148 -12170
rect 6089 -17990 6309 -12310
rect 11928 -17990 12148 -12310
rect 6089 -18130 12148 -17990
rect 12168 -12310 18227 -12170
rect 12168 -17990 12388 -12310
rect 18007 -17990 18227 -12310
rect 12168 -18130 18227 -17990
rect 18247 -12310 24306 -12170
rect 18247 -17990 18467 -12310
rect 18247 -18130 24306 -17990
rect -24306 -18370 -18247 -18230
rect -18467 -24190 -18247 -18370
rect -18227 -18370 -12168 -18230
rect -18227 -24190 -18007 -18370
rect -12388 -24190 -12168 -18370
rect -12148 -18370 -6089 -18230
rect -12148 -24190 -11928 -18370
rect -6309 -24190 -6089 -18370
rect -6069 -18370 -10 -18230
rect -6069 -24190 -5849 -18370
rect -230 -24190 -10 -18370
rect 10 -18370 6069 -18230
rect 10 -24190 230 -18370
rect 5849 -24190 6069 -18370
rect 6089 -18370 12148 -18230
rect 6089 -24190 6309 -18370
rect 11928 -24190 12148 -18370
rect 12168 -18370 18227 -18230
rect 12168 -24190 12388 -18370
rect 18007 -24190 18227 -18370
rect 18247 -18370 24306 -18230
rect 18247 -24190 18467 -18370
<< metal3 >>
rect -24306 24162 -18247 24190
rect -24306 18258 -18331 24162
rect -18267 18258 -18247 24162
rect -24306 18230 -18247 18258
rect -18227 24162 -12168 24190
rect -18227 18258 -12252 24162
rect -12188 18258 -12168 24162
rect -18227 18230 -12168 18258
rect -12148 24162 -6089 24190
rect -12148 18258 -6173 24162
rect -6109 18258 -6089 24162
rect -12148 18230 -6089 18258
rect -6069 24162 -10 24190
rect -6069 18258 -94 24162
rect -30 18258 -10 24162
rect -6069 18230 -10 18258
rect 10 24162 6069 24190
rect 10 18258 5985 24162
rect 6049 18258 6069 24162
rect 10 18230 6069 18258
rect 6089 24162 12148 24190
rect 6089 18258 12064 24162
rect 12128 18258 12148 24162
rect 6089 18230 12148 18258
rect 12168 24162 18227 24190
rect 12168 18258 18143 24162
rect 18207 18258 18227 24162
rect 12168 18230 18227 18258
rect 18247 24162 24306 24190
rect 18247 18258 24222 24162
rect 24286 18258 24306 24162
rect 18247 18230 24306 18258
rect -24306 18102 -18247 18130
rect -24306 12198 -18331 18102
rect -18267 12198 -18247 18102
rect -24306 12170 -18247 12198
rect -18227 18102 -12168 18130
rect -18227 12198 -12252 18102
rect -12188 12198 -12168 18102
rect -18227 12170 -12168 12198
rect -12148 18102 -6089 18130
rect -12148 12198 -6173 18102
rect -6109 12198 -6089 18102
rect -12148 12170 -6089 12198
rect -6069 18102 -10 18130
rect -6069 12198 -94 18102
rect -30 12198 -10 18102
rect -6069 12170 -10 12198
rect 10 18102 6069 18130
rect 10 12198 5985 18102
rect 6049 12198 6069 18102
rect 10 12170 6069 12198
rect 6089 18102 12148 18130
rect 6089 12198 12064 18102
rect 12128 12198 12148 18102
rect 6089 12170 12148 12198
rect 12168 18102 18227 18130
rect 12168 12198 18143 18102
rect 18207 12198 18227 18102
rect 12168 12170 18227 12198
rect 18247 18102 24306 18130
rect 18247 12198 24222 18102
rect 24286 12198 24306 18102
rect 18247 12170 24306 12198
rect -24306 12042 -18247 12070
rect -24306 6138 -18331 12042
rect -18267 6138 -18247 12042
rect -24306 6110 -18247 6138
rect -18227 12042 -12168 12070
rect -18227 6138 -12252 12042
rect -12188 6138 -12168 12042
rect -18227 6110 -12168 6138
rect -12148 12042 -6089 12070
rect -12148 6138 -6173 12042
rect -6109 6138 -6089 12042
rect -12148 6110 -6089 6138
rect -6069 12042 -10 12070
rect -6069 6138 -94 12042
rect -30 6138 -10 12042
rect -6069 6110 -10 6138
rect 10 12042 6069 12070
rect 10 6138 5985 12042
rect 6049 6138 6069 12042
rect 10 6110 6069 6138
rect 6089 12042 12148 12070
rect 6089 6138 12064 12042
rect 12128 6138 12148 12042
rect 6089 6110 12148 6138
rect 12168 12042 18227 12070
rect 12168 6138 18143 12042
rect 18207 6138 18227 12042
rect 12168 6110 18227 6138
rect 18247 12042 24306 12070
rect 18247 6138 24222 12042
rect 24286 6138 24306 12042
rect 18247 6110 24306 6138
rect -24306 5982 -18247 6010
rect -24306 78 -18331 5982
rect -18267 78 -18247 5982
rect -24306 50 -18247 78
rect -18227 5982 -12168 6010
rect -18227 78 -12252 5982
rect -12188 78 -12168 5982
rect -18227 50 -12168 78
rect -12148 5982 -6089 6010
rect -12148 78 -6173 5982
rect -6109 78 -6089 5982
rect -12148 50 -6089 78
rect -6069 5982 -10 6010
rect -6069 78 -94 5982
rect -30 78 -10 5982
rect -6069 50 -10 78
rect 10 5982 6069 6010
rect 10 78 5985 5982
rect 6049 78 6069 5982
rect 10 50 6069 78
rect 6089 5982 12148 6010
rect 6089 78 12064 5982
rect 12128 78 12148 5982
rect 6089 50 12148 78
rect 12168 5982 18227 6010
rect 12168 78 18143 5982
rect 18207 78 18227 5982
rect 12168 50 18227 78
rect 18247 5982 24306 6010
rect 18247 78 24222 5982
rect 24286 78 24306 5982
rect 18247 50 24306 78
rect -24306 -78 -18247 -50
rect -24306 -5982 -18331 -78
rect -18267 -5982 -18247 -78
rect -24306 -6010 -18247 -5982
rect -18227 -78 -12168 -50
rect -18227 -5982 -12252 -78
rect -12188 -5982 -12168 -78
rect -18227 -6010 -12168 -5982
rect -12148 -78 -6089 -50
rect -12148 -5982 -6173 -78
rect -6109 -5982 -6089 -78
rect -12148 -6010 -6089 -5982
rect -6069 -78 -10 -50
rect -6069 -5982 -94 -78
rect -30 -5982 -10 -78
rect -6069 -6010 -10 -5982
rect 10 -78 6069 -50
rect 10 -5982 5985 -78
rect 6049 -5982 6069 -78
rect 10 -6010 6069 -5982
rect 6089 -78 12148 -50
rect 6089 -5982 12064 -78
rect 12128 -5982 12148 -78
rect 6089 -6010 12148 -5982
rect 12168 -78 18227 -50
rect 12168 -5982 18143 -78
rect 18207 -5982 18227 -78
rect 12168 -6010 18227 -5982
rect 18247 -78 24306 -50
rect 18247 -5982 24222 -78
rect 24286 -5982 24306 -78
rect 18247 -6010 24306 -5982
rect -24306 -6138 -18247 -6110
rect -24306 -12042 -18331 -6138
rect -18267 -12042 -18247 -6138
rect -24306 -12070 -18247 -12042
rect -18227 -6138 -12168 -6110
rect -18227 -12042 -12252 -6138
rect -12188 -12042 -12168 -6138
rect -18227 -12070 -12168 -12042
rect -12148 -6138 -6089 -6110
rect -12148 -12042 -6173 -6138
rect -6109 -12042 -6089 -6138
rect -12148 -12070 -6089 -12042
rect -6069 -6138 -10 -6110
rect -6069 -12042 -94 -6138
rect -30 -12042 -10 -6138
rect -6069 -12070 -10 -12042
rect 10 -6138 6069 -6110
rect 10 -12042 5985 -6138
rect 6049 -12042 6069 -6138
rect 10 -12070 6069 -12042
rect 6089 -6138 12148 -6110
rect 6089 -12042 12064 -6138
rect 12128 -12042 12148 -6138
rect 6089 -12070 12148 -12042
rect 12168 -6138 18227 -6110
rect 12168 -12042 18143 -6138
rect 18207 -12042 18227 -6138
rect 12168 -12070 18227 -12042
rect 18247 -6138 24306 -6110
rect 18247 -12042 24222 -6138
rect 24286 -12042 24306 -6138
rect 18247 -12070 24306 -12042
rect -24306 -12198 -18247 -12170
rect -24306 -18102 -18331 -12198
rect -18267 -18102 -18247 -12198
rect -24306 -18130 -18247 -18102
rect -18227 -12198 -12168 -12170
rect -18227 -18102 -12252 -12198
rect -12188 -18102 -12168 -12198
rect -18227 -18130 -12168 -18102
rect -12148 -12198 -6089 -12170
rect -12148 -18102 -6173 -12198
rect -6109 -18102 -6089 -12198
rect -12148 -18130 -6089 -18102
rect -6069 -12198 -10 -12170
rect -6069 -18102 -94 -12198
rect -30 -18102 -10 -12198
rect -6069 -18130 -10 -18102
rect 10 -12198 6069 -12170
rect 10 -18102 5985 -12198
rect 6049 -18102 6069 -12198
rect 10 -18130 6069 -18102
rect 6089 -12198 12148 -12170
rect 6089 -18102 12064 -12198
rect 12128 -18102 12148 -12198
rect 6089 -18130 12148 -18102
rect 12168 -12198 18227 -12170
rect 12168 -18102 18143 -12198
rect 18207 -18102 18227 -12198
rect 12168 -18130 18227 -18102
rect 18247 -12198 24306 -12170
rect 18247 -18102 24222 -12198
rect 24286 -18102 24306 -12198
rect 18247 -18130 24306 -18102
rect -24306 -18258 -18247 -18230
rect -24306 -24162 -18331 -18258
rect -18267 -24162 -18247 -18258
rect -24306 -24190 -18247 -24162
rect -18227 -18258 -12168 -18230
rect -18227 -24162 -12252 -18258
rect -12188 -24162 -12168 -18258
rect -18227 -24190 -12168 -24162
rect -12148 -18258 -6089 -18230
rect -12148 -24162 -6173 -18258
rect -6109 -24162 -6089 -18258
rect -12148 -24190 -6089 -24162
rect -6069 -18258 -10 -18230
rect -6069 -24162 -94 -18258
rect -30 -24162 -10 -18258
rect -6069 -24190 -10 -24162
rect 10 -18258 6069 -18230
rect 10 -24162 5985 -18258
rect 6049 -24162 6069 -18258
rect 10 -24190 6069 -24162
rect 6089 -18258 12148 -18230
rect 6089 -24162 12064 -18258
rect 12128 -24162 12148 -18258
rect 6089 -24190 12148 -24162
rect 12168 -18258 18227 -18230
rect 12168 -24162 18143 -18258
rect 18207 -24162 18227 -18258
rect 12168 -24190 18227 -24162
rect 18247 -18258 24306 -18230
rect 18247 -24162 24222 -18258
rect 24286 -24162 24306 -18258
rect 18247 -24190 24306 -24162
<< via3 >>
rect -18331 18258 -18267 24162
rect -12252 18258 -12188 24162
rect -6173 18258 -6109 24162
rect -94 18258 -30 24162
rect 5985 18258 6049 24162
rect 12064 18258 12128 24162
rect 18143 18258 18207 24162
rect 24222 18258 24286 24162
rect -18331 12198 -18267 18102
rect -12252 12198 -12188 18102
rect -6173 12198 -6109 18102
rect -94 12198 -30 18102
rect 5985 12198 6049 18102
rect 12064 12198 12128 18102
rect 18143 12198 18207 18102
rect 24222 12198 24286 18102
rect -18331 6138 -18267 12042
rect -12252 6138 -12188 12042
rect -6173 6138 -6109 12042
rect -94 6138 -30 12042
rect 5985 6138 6049 12042
rect 12064 6138 12128 12042
rect 18143 6138 18207 12042
rect 24222 6138 24286 12042
rect -18331 78 -18267 5982
rect -12252 78 -12188 5982
rect -6173 78 -6109 5982
rect -94 78 -30 5982
rect 5985 78 6049 5982
rect 12064 78 12128 5982
rect 18143 78 18207 5982
rect 24222 78 24286 5982
rect -18331 -5982 -18267 -78
rect -12252 -5982 -12188 -78
rect -6173 -5982 -6109 -78
rect -94 -5982 -30 -78
rect 5985 -5982 6049 -78
rect 12064 -5982 12128 -78
rect 18143 -5982 18207 -78
rect 24222 -5982 24286 -78
rect -18331 -12042 -18267 -6138
rect -12252 -12042 -12188 -6138
rect -6173 -12042 -6109 -6138
rect -94 -12042 -30 -6138
rect 5985 -12042 6049 -6138
rect 12064 -12042 12128 -6138
rect 18143 -12042 18207 -6138
rect 24222 -12042 24286 -6138
rect -18331 -18102 -18267 -12198
rect -12252 -18102 -12188 -12198
rect -6173 -18102 -6109 -12198
rect -94 -18102 -30 -12198
rect 5985 -18102 6049 -12198
rect 12064 -18102 12128 -12198
rect 18143 -18102 18207 -12198
rect 24222 -18102 24286 -12198
rect -18331 -24162 -18267 -18258
rect -12252 -24162 -12188 -18258
rect -6173 -24162 -6109 -18258
rect -94 -24162 -30 -18258
rect 5985 -24162 6049 -18258
rect 12064 -24162 12128 -18258
rect 18143 -24162 18207 -18258
rect 24222 -24162 24286 -18258
<< mimcap >>
rect -24206 24050 -18446 24090
rect -24206 18370 -24166 24050
rect -18486 18370 -18446 24050
rect -24206 18330 -18446 18370
rect -18127 24050 -12367 24090
rect -18127 18370 -18087 24050
rect -12407 18370 -12367 24050
rect -18127 18330 -12367 18370
rect -12048 24050 -6288 24090
rect -12048 18370 -12008 24050
rect -6328 18370 -6288 24050
rect -12048 18330 -6288 18370
rect -5969 24050 -209 24090
rect -5969 18370 -5929 24050
rect -249 18370 -209 24050
rect -5969 18330 -209 18370
rect 110 24050 5870 24090
rect 110 18370 150 24050
rect 5830 18370 5870 24050
rect 110 18330 5870 18370
rect 6189 24050 11949 24090
rect 6189 18370 6229 24050
rect 11909 18370 11949 24050
rect 6189 18330 11949 18370
rect 12268 24050 18028 24090
rect 12268 18370 12308 24050
rect 17988 18370 18028 24050
rect 12268 18330 18028 18370
rect 18347 24050 24107 24090
rect 18347 18370 18387 24050
rect 24067 18370 24107 24050
rect 18347 18330 24107 18370
rect -24206 17990 -18446 18030
rect -24206 12310 -24166 17990
rect -18486 12310 -18446 17990
rect -24206 12270 -18446 12310
rect -18127 17990 -12367 18030
rect -18127 12310 -18087 17990
rect -12407 12310 -12367 17990
rect -18127 12270 -12367 12310
rect -12048 17990 -6288 18030
rect -12048 12310 -12008 17990
rect -6328 12310 -6288 17990
rect -12048 12270 -6288 12310
rect -5969 17990 -209 18030
rect -5969 12310 -5929 17990
rect -249 12310 -209 17990
rect -5969 12270 -209 12310
rect 110 17990 5870 18030
rect 110 12310 150 17990
rect 5830 12310 5870 17990
rect 110 12270 5870 12310
rect 6189 17990 11949 18030
rect 6189 12310 6229 17990
rect 11909 12310 11949 17990
rect 6189 12270 11949 12310
rect 12268 17990 18028 18030
rect 12268 12310 12308 17990
rect 17988 12310 18028 17990
rect 12268 12270 18028 12310
rect 18347 17990 24107 18030
rect 18347 12310 18387 17990
rect 24067 12310 24107 17990
rect 18347 12270 24107 12310
rect -24206 11930 -18446 11970
rect -24206 6250 -24166 11930
rect -18486 6250 -18446 11930
rect -24206 6210 -18446 6250
rect -18127 11930 -12367 11970
rect -18127 6250 -18087 11930
rect -12407 6250 -12367 11930
rect -18127 6210 -12367 6250
rect -12048 11930 -6288 11970
rect -12048 6250 -12008 11930
rect -6328 6250 -6288 11930
rect -12048 6210 -6288 6250
rect -5969 11930 -209 11970
rect -5969 6250 -5929 11930
rect -249 6250 -209 11930
rect -5969 6210 -209 6250
rect 110 11930 5870 11970
rect 110 6250 150 11930
rect 5830 6250 5870 11930
rect 110 6210 5870 6250
rect 6189 11930 11949 11970
rect 6189 6250 6229 11930
rect 11909 6250 11949 11930
rect 6189 6210 11949 6250
rect 12268 11930 18028 11970
rect 12268 6250 12308 11930
rect 17988 6250 18028 11930
rect 12268 6210 18028 6250
rect 18347 11930 24107 11970
rect 18347 6250 18387 11930
rect 24067 6250 24107 11930
rect 18347 6210 24107 6250
rect -24206 5870 -18446 5910
rect -24206 190 -24166 5870
rect -18486 190 -18446 5870
rect -24206 150 -18446 190
rect -18127 5870 -12367 5910
rect -18127 190 -18087 5870
rect -12407 190 -12367 5870
rect -18127 150 -12367 190
rect -12048 5870 -6288 5910
rect -12048 190 -12008 5870
rect -6328 190 -6288 5870
rect -12048 150 -6288 190
rect -5969 5870 -209 5910
rect -5969 190 -5929 5870
rect -249 190 -209 5870
rect -5969 150 -209 190
rect 110 5870 5870 5910
rect 110 190 150 5870
rect 5830 190 5870 5870
rect 110 150 5870 190
rect 6189 5870 11949 5910
rect 6189 190 6229 5870
rect 11909 190 11949 5870
rect 6189 150 11949 190
rect 12268 5870 18028 5910
rect 12268 190 12308 5870
rect 17988 190 18028 5870
rect 12268 150 18028 190
rect 18347 5870 24107 5910
rect 18347 190 18387 5870
rect 24067 190 24107 5870
rect 18347 150 24107 190
rect -24206 -190 -18446 -150
rect -24206 -5870 -24166 -190
rect -18486 -5870 -18446 -190
rect -24206 -5910 -18446 -5870
rect -18127 -190 -12367 -150
rect -18127 -5870 -18087 -190
rect -12407 -5870 -12367 -190
rect -18127 -5910 -12367 -5870
rect -12048 -190 -6288 -150
rect -12048 -5870 -12008 -190
rect -6328 -5870 -6288 -190
rect -12048 -5910 -6288 -5870
rect -5969 -190 -209 -150
rect -5969 -5870 -5929 -190
rect -249 -5870 -209 -190
rect -5969 -5910 -209 -5870
rect 110 -190 5870 -150
rect 110 -5870 150 -190
rect 5830 -5870 5870 -190
rect 110 -5910 5870 -5870
rect 6189 -190 11949 -150
rect 6189 -5870 6229 -190
rect 11909 -5870 11949 -190
rect 6189 -5910 11949 -5870
rect 12268 -190 18028 -150
rect 12268 -5870 12308 -190
rect 17988 -5870 18028 -190
rect 12268 -5910 18028 -5870
rect 18347 -190 24107 -150
rect 18347 -5870 18387 -190
rect 24067 -5870 24107 -190
rect 18347 -5910 24107 -5870
rect -24206 -6250 -18446 -6210
rect -24206 -11930 -24166 -6250
rect -18486 -11930 -18446 -6250
rect -24206 -11970 -18446 -11930
rect -18127 -6250 -12367 -6210
rect -18127 -11930 -18087 -6250
rect -12407 -11930 -12367 -6250
rect -18127 -11970 -12367 -11930
rect -12048 -6250 -6288 -6210
rect -12048 -11930 -12008 -6250
rect -6328 -11930 -6288 -6250
rect -12048 -11970 -6288 -11930
rect -5969 -6250 -209 -6210
rect -5969 -11930 -5929 -6250
rect -249 -11930 -209 -6250
rect -5969 -11970 -209 -11930
rect 110 -6250 5870 -6210
rect 110 -11930 150 -6250
rect 5830 -11930 5870 -6250
rect 110 -11970 5870 -11930
rect 6189 -6250 11949 -6210
rect 6189 -11930 6229 -6250
rect 11909 -11930 11949 -6250
rect 6189 -11970 11949 -11930
rect 12268 -6250 18028 -6210
rect 12268 -11930 12308 -6250
rect 17988 -11930 18028 -6250
rect 12268 -11970 18028 -11930
rect 18347 -6250 24107 -6210
rect 18347 -11930 18387 -6250
rect 24067 -11930 24107 -6250
rect 18347 -11970 24107 -11930
rect -24206 -12310 -18446 -12270
rect -24206 -17990 -24166 -12310
rect -18486 -17990 -18446 -12310
rect -24206 -18030 -18446 -17990
rect -18127 -12310 -12367 -12270
rect -18127 -17990 -18087 -12310
rect -12407 -17990 -12367 -12310
rect -18127 -18030 -12367 -17990
rect -12048 -12310 -6288 -12270
rect -12048 -17990 -12008 -12310
rect -6328 -17990 -6288 -12310
rect -12048 -18030 -6288 -17990
rect -5969 -12310 -209 -12270
rect -5969 -17990 -5929 -12310
rect -249 -17990 -209 -12310
rect -5969 -18030 -209 -17990
rect 110 -12310 5870 -12270
rect 110 -17990 150 -12310
rect 5830 -17990 5870 -12310
rect 110 -18030 5870 -17990
rect 6189 -12310 11949 -12270
rect 6189 -17990 6229 -12310
rect 11909 -17990 11949 -12310
rect 6189 -18030 11949 -17990
rect 12268 -12310 18028 -12270
rect 12268 -17990 12308 -12310
rect 17988 -17990 18028 -12310
rect 12268 -18030 18028 -17990
rect 18347 -12310 24107 -12270
rect 18347 -17990 18387 -12310
rect 24067 -17990 24107 -12310
rect 18347 -18030 24107 -17990
rect -24206 -18370 -18446 -18330
rect -24206 -24050 -24166 -18370
rect -18486 -24050 -18446 -18370
rect -24206 -24090 -18446 -24050
rect -18127 -18370 -12367 -18330
rect -18127 -24050 -18087 -18370
rect -12407 -24050 -12367 -18370
rect -18127 -24090 -12367 -24050
rect -12048 -18370 -6288 -18330
rect -12048 -24050 -12008 -18370
rect -6328 -24050 -6288 -18370
rect -12048 -24090 -6288 -24050
rect -5969 -18370 -209 -18330
rect -5969 -24050 -5929 -18370
rect -249 -24050 -209 -18370
rect -5969 -24090 -209 -24050
rect 110 -18370 5870 -18330
rect 110 -24050 150 -18370
rect 5830 -24050 5870 -18370
rect 110 -24090 5870 -24050
rect 6189 -18370 11949 -18330
rect 6189 -24050 6229 -18370
rect 11909 -24050 11949 -18370
rect 6189 -24090 11949 -24050
rect 12268 -18370 18028 -18330
rect 12268 -24050 12308 -18370
rect 17988 -24050 18028 -18370
rect 12268 -24090 18028 -24050
rect 18347 -18370 24107 -18330
rect 18347 -24050 18387 -18370
rect 24067 -24050 24107 -18370
rect 18347 -24090 24107 -24050
<< mimcapcontact >>
rect -24166 18370 -18486 24050
rect -18087 18370 -12407 24050
rect -12008 18370 -6328 24050
rect -5929 18370 -249 24050
rect 150 18370 5830 24050
rect 6229 18370 11909 24050
rect 12308 18370 17988 24050
rect 18387 18370 24067 24050
rect -24166 12310 -18486 17990
rect -18087 12310 -12407 17990
rect -12008 12310 -6328 17990
rect -5929 12310 -249 17990
rect 150 12310 5830 17990
rect 6229 12310 11909 17990
rect 12308 12310 17988 17990
rect 18387 12310 24067 17990
rect -24166 6250 -18486 11930
rect -18087 6250 -12407 11930
rect -12008 6250 -6328 11930
rect -5929 6250 -249 11930
rect 150 6250 5830 11930
rect 6229 6250 11909 11930
rect 12308 6250 17988 11930
rect 18387 6250 24067 11930
rect -24166 190 -18486 5870
rect -18087 190 -12407 5870
rect -12008 190 -6328 5870
rect -5929 190 -249 5870
rect 150 190 5830 5870
rect 6229 190 11909 5870
rect 12308 190 17988 5870
rect 18387 190 24067 5870
rect -24166 -5870 -18486 -190
rect -18087 -5870 -12407 -190
rect -12008 -5870 -6328 -190
rect -5929 -5870 -249 -190
rect 150 -5870 5830 -190
rect 6229 -5870 11909 -190
rect 12308 -5870 17988 -190
rect 18387 -5870 24067 -190
rect -24166 -11930 -18486 -6250
rect -18087 -11930 -12407 -6250
rect -12008 -11930 -6328 -6250
rect -5929 -11930 -249 -6250
rect 150 -11930 5830 -6250
rect 6229 -11930 11909 -6250
rect 12308 -11930 17988 -6250
rect 18387 -11930 24067 -6250
rect -24166 -17990 -18486 -12310
rect -18087 -17990 -12407 -12310
rect -12008 -17990 -6328 -12310
rect -5929 -17990 -249 -12310
rect 150 -17990 5830 -12310
rect 6229 -17990 11909 -12310
rect 12308 -17990 17988 -12310
rect 18387 -17990 24067 -12310
rect -24166 -24050 -18486 -18370
rect -18087 -24050 -12407 -18370
rect -12008 -24050 -6328 -18370
rect -5929 -24050 -249 -18370
rect 150 -24050 5830 -18370
rect 6229 -24050 11909 -18370
rect 12308 -24050 17988 -18370
rect 18387 -24050 24067 -18370
<< metal4 >>
rect -21378 24051 -21274 24240
rect -18378 24178 -18274 24240
rect -18378 24162 -18251 24178
rect -24167 24050 -18485 24051
rect -24167 18370 -24166 24050
rect -18486 18370 -18485 24050
rect -24167 18369 -18485 18370
rect -21378 17991 -21274 18369
rect -18378 18258 -18331 24162
rect -18267 18258 -18251 24162
rect -15299 24051 -15195 24240
rect -12299 24178 -12195 24240
rect -12299 24162 -12172 24178
rect -18088 24050 -12406 24051
rect -18088 18370 -18087 24050
rect -12407 18370 -12406 24050
rect -18088 18369 -12406 18370
rect -18378 18242 -18251 18258
rect -18378 18118 -18274 18242
rect -18378 18102 -18251 18118
rect -24167 17990 -18485 17991
rect -24167 12310 -24166 17990
rect -18486 12310 -18485 17990
rect -24167 12309 -18485 12310
rect -21378 11931 -21274 12309
rect -18378 12198 -18331 18102
rect -18267 12198 -18251 18102
rect -15299 17991 -15195 18369
rect -12299 18258 -12252 24162
rect -12188 18258 -12172 24162
rect -9220 24051 -9116 24240
rect -6220 24178 -6116 24240
rect -6220 24162 -6093 24178
rect -12009 24050 -6327 24051
rect -12009 18370 -12008 24050
rect -6328 18370 -6327 24050
rect -12009 18369 -6327 18370
rect -12299 18242 -12172 18258
rect -12299 18118 -12195 18242
rect -12299 18102 -12172 18118
rect -18088 17990 -12406 17991
rect -18088 12310 -18087 17990
rect -12407 12310 -12406 17990
rect -18088 12309 -12406 12310
rect -18378 12182 -18251 12198
rect -18378 12058 -18274 12182
rect -18378 12042 -18251 12058
rect -24167 11930 -18485 11931
rect -24167 6250 -24166 11930
rect -18486 6250 -18485 11930
rect -24167 6249 -18485 6250
rect -21378 5871 -21274 6249
rect -18378 6138 -18331 12042
rect -18267 6138 -18251 12042
rect -15299 11931 -15195 12309
rect -12299 12198 -12252 18102
rect -12188 12198 -12172 18102
rect -9220 17991 -9116 18369
rect -6220 18258 -6173 24162
rect -6109 18258 -6093 24162
rect -3141 24051 -3037 24240
rect -141 24178 -37 24240
rect -141 24162 -14 24178
rect -5930 24050 -248 24051
rect -5930 18370 -5929 24050
rect -249 18370 -248 24050
rect -5930 18369 -248 18370
rect -6220 18242 -6093 18258
rect -6220 18118 -6116 18242
rect -6220 18102 -6093 18118
rect -12009 17990 -6327 17991
rect -12009 12310 -12008 17990
rect -6328 12310 -6327 17990
rect -12009 12309 -6327 12310
rect -12299 12182 -12172 12198
rect -12299 12058 -12195 12182
rect -12299 12042 -12172 12058
rect -18088 11930 -12406 11931
rect -18088 6250 -18087 11930
rect -12407 6250 -12406 11930
rect -18088 6249 -12406 6250
rect -18378 6122 -18251 6138
rect -18378 5998 -18274 6122
rect -18378 5982 -18251 5998
rect -24167 5870 -18485 5871
rect -24167 190 -24166 5870
rect -18486 190 -18485 5870
rect -24167 189 -18485 190
rect -21378 -189 -21274 189
rect -18378 78 -18331 5982
rect -18267 78 -18251 5982
rect -15299 5871 -15195 6249
rect -12299 6138 -12252 12042
rect -12188 6138 -12172 12042
rect -9220 11931 -9116 12309
rect -6220 12198 -6173 18102
rect -6109 12198 -6093 18102
rect -3141 17991 -3037 18369
rect -141 18258 -94 24162
rect -30 18258 -14 24162
rect 2938 24051 3042 24240
rect 5938 24178 6042 24240
rect 5938 24162 6065 24178
rect 149 24050 5831 24051
rect 149 18370 150 24050
rect 5830 18370 5831 24050
rect 149 18369 5831 18370
rect -141 18242 -14 18258
rect -141 18118 -37 18242
rect -141 18102 -14 18118
rect -5930 17990 -248 17991
rect -5930 12310 -5929 17990
rect -249 12310 -248 17990
rect -5930 12309 -248 12310
rect -6220 12182 -6093 12198
rect -6220 12058 -6116 12182
rect -6220 12042 -6093 12058
rect -12009 11930 -6327 11931
rect -12009 6250 -12008 11930
rect -6328 6250 -6327 11930
rect -12009 6249 -6327 6250
rect -12299 6122 -12172 6138
rect -12299 5998 -12195 6122
rect -12299 5982 -12172 5998
rect -18088 5870 -12406 5871
rect -18088 190 -18087 5870
rect -12407 190 -12406 5870
rect -18088 189 -12406 190
rect -18378 62 -18251 78
rect -18378 -62 -18274 62
rect -18378 -78 -18251 -62
rect -24167 -190 -18485 -189
rect -24167 -5870 -24166 -190
rect -18486 -5870 -18485 -190
rect -24167 -5871 -18485 -5870
rect -21378 -6249 -21274 -5871
rect -18378 -5982 -18331 -78
rect -18267 -5982 -18251 -78
rect -15299 -189 -15195 189
rect -12299 78 -12252 5982
rect -12188 78 -12172 5982
rect -9220 5871 -9116 6249
rect -6220 6138 -6173 12042
rect -6109 6138 -6093 12042
rect -3141 11931 -3037 12309
rect -141 12198 -94 18102
rect -30 12198 -14 18102
rect 2938 17991 3042 18369
rect 5938 18258 5985 24162
rect 6049 18258 6065 24162
rect 9017 24051 9121 24240
rect 12017 24178 12121 24240
rect 12017 24162 12144 24178
rect 6228 24050 11910 24051
rect 6228 18370 6229 24050
rect 11909 18370 11910 24050
rect 6228 18369 11910 18370
rect 5938 18242 6065 18258
rect 5938 18118 6042 18242
rect 5938 18102 6065 18118
rect 149 17990 5831 17991
rect 149 12310 150 17990
rect 5830 12310 5831 17990
rect 149 12309 5831 12310
rect -141 12182 -14 12198
rect -141 12058 -37 12182
rect -141 12042 -14 12058
rect -5930 11930 -248 11931
rect -5930 6250 -5929 11930
rect -249 6250 -248 11930
rect -5930 6249 -248 6250
rect -6220 6122 -6093 6138
rect -6220 5998 -6116 6122
rect -6220 5982 -6093 5998
rect -12009 5870 -6327 5871
rect -12009 190 -12008 5870
rect -6328 190 -6327 5870
rect -12009 189 -6327 190
rect -12299 62 -12172 78
rect -12299 -62 -12195 62
rect -12299 -78 -12172 -62
rect -18088 -190 -12406 -189
rect -18088 -5870 -18087 -190
rect -12407 -5870 -12406 -190
rect -18088 -5871 -12406 -5870
rect -18378 -5998 -18251 -5982
rect -18378 -6122 -18274 -5998
rect -18378 -6138 -18251 -6122
rect -24167 -6250 -18485 -6249
rect -24167 -11930 -24166 -6250
rect -18486 -11930 -18485 -6250
rect -24167 -11931 -18485 -11930
rect -21378 -12309 -21274 -11931
rect -18378 -12042 -18331 -6138
rect -18267 -12042 -18251 -6138
rect -15299 -6249 -15195 -5871
rect -12299 -5982 -12252 -78
rect -12188 -5982 -12172 -78
rect -9220 -189 -9116 189
rect -6220 78 -6173 5982
rect -6109 78 -6093 5982
rect -3141 5871 -3037 6249
rect -141 6138 -94 12042
rect -30 6138 -14 12042
rect 2938 11931 3042 12309
rect 5938 12198 5985 18102
rect 6049 12198 6065 18102
rect 9017 17991 9121 18369
rect 12017 18258 12064 24162
rect 12128 18258 12144 24162
rect 15096 24051 15200 24240
rect 18096 24178 18200 24240
rect 18096 24162 18223 24178
rect 12307 24050 17989 24051
rect 12307 18370 12308 24050
rect 17988 18370 17989 24050
rect 12307 18369 17989 18370
rect 12017 18242 12144 18258
rect 12017 18118 12121 18242
rect 12017 18102 12144 18118
rect 6228 17990 11910 17991
rect 6228 12310 6229 17990
rect 11909 12310 11910 17990
rect 6228 12309 11910 12310
rect 5938 12182 6065 12198
rect 5938 12058 6042 12182
rect 5938 12042 6065 12058
rect 149 11930 5831 11931
rect 149 6250 150 11930
rect 5830 6250 5831 11930
rect 149 6249 5831 6250
rect -141 6122 -14 6138
rect -141 5998 -37 6122
rect -141 5982 -14 5998
rect -5930 5870 -248 5871
rect -5930 190 -5929 5870
rect -249 190 -248 5870
rect -5930 189 -248 190
rect -6220 62 -6093 78
rect -6220 -62 -6116 62
rect -6220 -78 -6093 -62
rect -12009 -190 -6327 -189
rect -12009 -5870 -12008 -190
rect -6328 -5870 -6327 -190
rect -12009 -5871 -6327 -5870
rect -12299 -5998 -12172 -5982
rect -12299 -6122 -12195 -5998
rect -12299 -6138 -12172 -6122
rect -18088 -6250 -12406 -6249
rect -18088 -11930 -18087 -6250
rect -12407 -11930 -12406 -6250
rect -18088 -11931 -12406 -11930
rect -18378 -12058 -18251 -12042
rect -18378 -12182 -18274 -12058
rect -18378 -12198 -18251 -12182
rect -24167 -12310 -18485 -12309
rect -24167 -17990 -24166 -12310
rect -18486 -17990 -18485 -12310
rect -24167 -17991 -18485 -17990
rect -21378 -18369 -21274 -17991
rect -18378 -18102 -18331 -12198
rect -18267 -18102 -18251 -12198
rect -15299 -12309 -15195 -11931
rect -12299 -12042 -12252 -6138
rect -12188 -12042 -12172 -6138
rect -9220 -6249 -9116 -5871
rect -6220 -5982 -6173 -78
rect -6109 -5982 -6093 -78
rect -3141 -189 -3037 189
rect -141 78 -94 5982
rect -30 78 -14 5982
rect 2938 5871 3042 6249
rect 5938 6138 5985 12042
rect 6049 6138 6065 12042
rect 9017 11931 9121 12309
rect 12017 12198 12064 18102
rect 12128 12198 12144 18102
rect 15096 17991 15200 18369
rect 18096 18258 18143 24162
rect 18207 18258 18223 24162
rect 21175 24051 21279 24240
rect 24175 24178 24279 24240
rect 24175 24162 24302 24178
rect 18386 24050 24068 24051
rect 18386 18370 18387 24050
rect 24067 18370 24068 24050
rect 18386 18369 24068 18370
rect 18096 18242 18223 18258
rect 18096 18118 18200 18242
rect 18096 18102 18223 18118
rect 12307 17990 17989 17991
rect 12307 12310 12308 17990
rect 17988 12310 17989 17990
rect 12307 12309 17989 12310
rect 12017 12182 12144 12198
rect 12017 12058 12121 12182
rect 12017 12042 12144 12058
rect 6228 11930 11910 11931
rect 6228 6250 6229 11930
rect 11909 6250 11910 11930
rect 6228 6249 11910 6250
rect 5938 6122 6065 6138
rect 5938 5998 6042 6122
rect 5938 5982 6065 5998
rect 149 5870 5831 5871
rect 149 190 150 5870
rect 5830 190 5831 5870
rect 149 189 5831 190
rect -141 62 -14 78
rect -141 -62 -37 62
rect -141 -78 -14 -62
rect -5930 -190 -248 -189
rect -5930 -5870 -5929 -190
rect -249 -5870 -248 -190
rect -5930 -5871 -248 -5870
rect -6220 -5998 -6093 -5982
rect -6220 -6122 -6116 -5998
rect -6220 -6138 -6093 -6122
rect -12009 -6250 -6327 -6249
rect -12009 -11930 -12008 -6250
rect -6328 -11930 -6327 -6250
rect -12009 -11931 -6327 -11930
rect -12299 -12058 -12172 -12042
rect -12299 -12182 -12195 -12058
rect -12299 -12198 -12172 -12182
rect -18088 -12310 -12406 -12309
rect -18088 -17990 -18087 -12310
rect -12407 -17990 -12406 -12310
rect -18088 -17991 -12406 -17990
rect -18378 -18118 -18251 -18102
rect -18378 -18242 -18274 -18118
rect -18378 -18258 -18251 -18242
rect -24167 -18370 -18485 -18369
rect -24167 -24050 -24166 -18370
rect -18486 -24050 -18485 -18370
rect -24167 -24051 -18485 -24050
rect -21378 -24240 -21274 -24051
rect -18378 -24162 -18331 -18258
rect -18267 -24162 -18251 -18258
rect -15299 -18369 -15195 -17991
rect -12299 -18102 -12252 -12198
rect -12188 -18102 -12172 -12198
rect -9220 -12309 -9116 -11931
rect -6220 -12042 -6173 -6138
rect -6109 -12042 -6093 -6138
rect -3141 -6249 -3037 -5871
rect -141 -5982 -94 -78
rect -30 -5982 -14 -78
rect 2938 -189 3042 189
rect 5938 78 5985 5982
rect 6049 78 6065 5982
rect 9017 5871 9121 6249
rect 12017 6138 12064 12042
rect 12128 6138 12144 12042
rect 15096 11931 15200 12309
rect 18096 12198 18143 18102
rect 18207 12198 18223 18102
rect 21175 17991 21279 18369
rect 24175 18258 24222 24162
rect 24286 18258 24302 24162
rect 24175 18242 24302 18258
rect 24175 18118 24279 18242
rect 24175 18102 24302 18118
rect 18386 17990 24068 17991
rect 18386 12310 18387 17990
rect 24067 12310 24068 17990
rect 18386 12309 24068 12310
rect 18096 12182 18223 12198
rect 18096 12058 18200 12182
rect 18096 12042 18223 12058
rect 12307 11930 17989 11931
rect 12307 6250 12308 11930
rect 17988 6250 17989 11930
rect 12307 6249 17989 6250
rect 12017 6122 12144 6138
rect 12017 5998 12121 6122
rect 12017 5982 12144 5998
rect 6228 5870 11910 5871
rect 6228 190 6229 5870
rect 11909 190 11910 5870
rect 6228 189 11910 190
rect 5938 62 6065 78
rect 5938 -62 6042 62
rect 5938 -78 6065 -62
rect 149 -190 5831 -189
rect 149 -5870 150 -190
rect 5830 -5870 5831 -190
rect 149 -5871 5831 -5870
rect -141 -5998 -14 -5982
rect -141 -6122 -37 -5998
rect -141 -6138 -14 -6122
rect -5930 -6250 -248 -6249
rect -5930 -11930 -5929 -6250
rect -249 -11930 -248 -6250
rect -5930 -11931 -248 -11930
rect -6220 -12058 -6093 -12042
rect -6220 -12182 -6116 -12058
rect -6220 -12198 -6093 -12182
rect -12009 -12310 -6327 -12309
rect -12009 -17990 -12008 -12310
rect -6328 -17990 -6327 -12310
rect -12009 -17991 -6327 -17990
rect -12299 -18118 -12172 -18102
rect -12299 -18242 -12195 -18118
rect -12299 -18258 -12172 -18242
rect -18088 -18370 -12406 -18369
rect -18088 -24050 -18087 -18370
rect -12407 -24050 -12406 -18370
rect -18088 -24051 -12406 -24050
rect -18378 -24178 -18251 -24162
rect -18378 -24240 -18274 -24178
rect -15299 -24240 -15195 -24051
rect -12299 -24162 -12252 -18258
rect -12188 -24162 -12172 -18258
rect -9220 -18369 -9116 -17991
rect -6220 -18102 -6173 -12198
rect -6109 -18102 -6093 -12198
rect -3141 -12309 -3037 -11931
rect -141 -12042 -94 -6138
rect -30 -12042 -14 -6138
rect 2938 -6249 3042 -5871
rect 5938 -5982 5985 -78
rect 6049 -5982 6065 -78
rect 9017 -189 9121 189
rect 12017 78 12064 5982
rect 12128 78 12144 5982
rect 15096 5871 15200 6249
rect 18096 6138 18143 12042
rect 18207 6138 18223 12042
rect 21175 11931 21279 12309
rect 24175 12198 24222 18102
rect 24286 12198 24302 18102
rect 24175 12182 24302 12198
rect 24175 12058 24279 12182
rect 24175 12042 24302 12058
rect 18386 11930 24068 11931
rect 18386 6250 18387 11930
rect 24067 6250 24068 11930
rect 18386 6249 24068 6250
rect 18096 6122 18223 6138
rect 18096 5998 18200 6122
rect 18096 5982 18223 5998
rect 12307 5870 17989 5871
rect 12307 190 12308 5870
rect 17988 190 17989 5870
rect 12307 189 17989 190
rect 12017 62 12144 78
rect 12017 -62 12121 62
rect 12017 -78 12144 -62
rect 6228 -190 11910 -189
rect 6228 -5870 6229 -190
rect 11909 -5870 11910 -190
rect 6228 -5871 11910 -5870
rect 5938 -5998 6065 -5982
rect 5938 -6122 6042 -5998
rect 5938 -6138 6065 -6122
rect 149 -6250 5831 -6249
rect 149 -11930 150 -6250
rect 5830 -11930 5831 -6250
rect 149 -11931 5831 -11930
rect -141 -12058 -14 -12042
rect -141 -12182 -37 -12058
rect -141 -12198 -14 -12182
rect -5930 -12310 -248 -12309
rect -5930 -17990 -5929 -12310
rect -249 -17990 -248 -12310
rect -5930 -17991 -248 -17990
rect -6220 -18118 -6093 -18102
rect -6220 -18242 -6116 -18118
rect -6220 -18258 -6093 -18242
rect -12009 -18370 -6327 -18369
rect -12009 -24050 -12008 -18370
rect -6328 -24050 -6327 -18370
rect -12009 -24051 -6327 -24050
rect -12299 -24178 -12172 -24162
rect -12299 -24240 -12195 -24178
rect -9220 -24240 -9116 -24051
rect -6220 -24162 -6173 -18258
rect -6109 -24162 -6093 -18258
rect -3141 -18369 -3037 -17991
rect -141 -18102 -94 -12198
rect -30 -18102 -14 -12198
rect 2938 -12309 3042 -11931
rect 5938 -12042 5985 -6138
rect 6049 -12042 6065 -6138
rect 9017 -6249 9121 -5871
rect 12017 -5982 12064 -78
rect 12128 -5982 12144 -78
rect 15096 -189 15200 189
rect 18096 78 18143 5982
rect 18207 78 18223 5982
rect 21175 5871 21279 6249
rect 24175 6138 24222 12042
rect 24286 6138 24302 12042
rect 24175 6122 24302 6138
rect 24175 5998 24279 6122
rect 24175 5982 24302 5998
rect 18386 5870 24068 5871
rect 18386 190 18387 5870
rect 24067 190 24068 5870
rect 18386 189 24068 190
rect 18096 62 18223 78
rect 18096 -62 18200 62
rect 18096 -78 18223 -62
rect 12307 -190 17989 -189
rect 12307 -5870 12308 -190
rect 17988 -5870 17989 -190
rect 12307 -5871 17989 -5870
rect 12017 -5998 12144 -5982
rect 12017 -6122 12121 -5998
rect 12017 -6138 12144 -6122
rect 6228 -6250 11910 -6249
rect 6228 -11930 6229 -6250
rect 11909 -11930 11910 -6250
rect 6228 -11931 11910 -11930
rect 5938 -12058 6065 -12042
rect 5938 -12182 6042 -12058
rect 5938 -12198 6065 -12182
rect 149 -12310 5831 -12309
rect 149 -17990 150 -12310
rect 5830 -17990 5831 -12310
rect 149 -17991 5831 -17990
rect -141 -18118 -14 -18102
rect -141 -18242 -37 -18118
rect -141 -18258 -14 -18242
rect -5930 -18370 -248 -18369
rect -5930 -24050 -5929 -18370
rect -249 -24050 -248 -18370
rect -5930 -24051 -248 -24050
rect -6220 -24178 -6093 -24162
rect -6220 -24240 -6116 -24178
rect -3141 -24240 -3037 -24051
rect -141 -24162 -94 -18258
rect -30 -24162 -14 -18258
rect 2938 -18369 3042 -17991
rect 5938 -18102 5985 -12198
rect 6049 -18102 6065 -12198
rect 9017 -12309 9121 -11931
rect 12017 -12042 12064 -6138
rect 12128 -12042 12144 -6138
rect 15096 -6249 15200 -5871
rect 18096 -5982 18143 -78
rect 18207 -5982 18223 -78
rect 21175 -189 21279 189
rect 24175 78 24222 5982
rect 24286 78 24302 5982
rect 24175 62 24302 78
rect 24175 -62 24279 62
rect 24175 -78 24302 -62
rect 18386 -190 24068 -189
rect 18386 -5870 18387 -190
rect 24067 -5870 24068 -190
rect 18386 -5871 24068 -5870
rect 18096 -5998 18223 -5982
rect 18096 -6122 18200 -5998
rect 18096 -6138 18223 -6122
rect 12307 -6250 17989 -6249
rect 12307 -11930 12308 -6250
rect 17988 -11930 17989 -6250
rect 12307 -11931 17989 -11930
rect 12017 -12058 12144 -12042
rect 12017 -12182 12121 -12058
rect 12017 -12198 12144 -12182
rect 6228 -12310 11910 -12309
rect 6228 -17990 6229 -12310
rect 11909 -17990 11910 -12310
rect 6228 -17991 11910 -17990
rect 5938 -18118 6065 -18102
rect 5938 -18242 6042 -18118
rect 5938 -18258 6065 -18242
rect 149 -18370 5831 -18369
rect 149 -24050 150 -18370
rect 5830 -24050 5831 -18370
rect 149 -24051 5831 -24050
rect -141 -24178 -14 -24162
rect -141 -24240 -37 -24178
rect 2938 -24240 3042 -24051
rect 5938 -24162 5985 -18258
rect 6049 -24162 6065 -18258
rect 9017 -18369 9121 -17991
rect 12017 -18102 12064 -12198
rect 12128 -18102 12144 -12198
rect 15096 -12309 15200 -11931
rect 18096 -12042 18143 -6138
rect 18207 -12042 18223 -6138
rect 21175 -6249 21279 -5871
rect 24175 -5982 24222 -78
rect 24286 -5982 24302 -78
rect 24175 -5998 24302 -5982
rect 24175 -6122 24279 -5998
rect 24175 -6138 24302 -6122
rect 18386 -6250 24068 -6249
rect 18386 -11930 18387 -6250
rect 24067 -11930 24068 -6250
rect 18386 -11931 24068 -11930
rect 18096 -12058 18223 -12042
rect 18096 -12182 18200 -12058
rect 18096 -12198 18223 -12182
rect 12307 -12310 17989 -12309
rect 12307 -17990 12308 -12310
rect 17988 -17990 17989 -12310
rect 12307 -17991 17989 -17990
rect 12017 -18118 12144 -18102
rect 12017 -18242 12121 -18118
rect 12017 -18258 12144 -18242
rect 6228 -18370 11910 -18369
rect 6228 -24050 6229 -18370
rect 11909 -24050 11910 -18370
rect 6228 -24051 11910 -24050
rect 5938 -24178 6065 -24162
rect 5938 -24240 6042 -24178
rect 9017 -24240 9121 -24051
rect 12017 -24162 12064 -18258
rect 12128 -24162 12144 -18258
rect 15096 -18369 15200 -17991
rect 18096 -18102 18143 -12198
rect 18207 -18102 18223 -12198
rect 21175 -12309 21279 -11931
rect 24175 -12042 24222 -6138
rect 24286 -12042 24302 -6138
rect 24175 -12058 24302 -12042
rect 24175 -12182 24279 -12058
rect 24175 -12198 24302 -12182
rect 18386 -12310 24068 -12309
rect 18386 -17990 18387 -12310
rect 24067 -17990 24068 -12310
rect 18386 -17991 24068 -17990
rect 18096 -18118 18223 -18102
rect 18096 -18242 18200 -18118
rect 18096 -18258 18223 -18242
rect 12307 -18370 17989 -18369
rect 12307 -24050 12308 -18370
rect 17988 -24050 17989 -18370
rect 12307 -24051 17989 -24050
rect 12017 -24178 12144 -24162
rect 12017 -24240 12121 -24178
rect 15096 -24240 15200 -24051
rect 18096 -24162 18143 -18258
rect 18207 -24162 18223 -18258
rect 21175 -18369 21279 -17991
rect 24175 -18102 24222 -12198
rect 24286 -18102 24302 -12198
rect 24175 -18118 24302 -18102
rect 24175 -18242 24279 -18118
rect 24175 -18258 24302 -18242
rect 18386 -18370 24068 -18369
rect 18386 -24050 18387 -18370
rect 24067 -24050 24068 -18370
rect 18386 -24051 24068 -24050
rect 18096 -24178 18223 -24162
rect 18096 -24240 18200 -24178
rect 21175 -24240 21279 -24051
rect 24175 -24162 24222 -18258
rect 24286 -24162 24302 -18258
rect 24175 -24178 24302 -24162
rect 24175 -24240 24279 -24178
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX 18247 18230 24207 24190
string parameters w 28.8 l 28.8 val 1.68k carea 2.00 cperi 0.19 nx 8 ny 8 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
string library sky130
<< end >>
