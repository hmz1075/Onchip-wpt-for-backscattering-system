* NGSPICE file created from FINAL_without_ind.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_lvt_4QC8GG a_n93_n5000# w_n231_n5219# a_n35_n5097#
+ a_35_n5000# VSUBS
X0 a_35_n5000# a_n35_n5097# a_n93_n5000# w_n231_n5219# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+07u l=350000u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_8K7EBA w_n231_n2210# a_n93_n2000# a_35_n2000#
+ a_n35_n2088#
X0 a_35_n2000# a_n35_n2088# a_n93_n2000# w_n231_n2210# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+07u l=350000u
.ends

.subckt Comparator_jafar VSS VIN- VINp VOUT
Xsky130_fd_pr__pfet_01v8_lvt_4QC8GG_0 VIN- VIN- a_3872_2262# m1_7222_1296# VSS sky130_fd_pr__pfet_01v8_lvt_4QC8GG
Xsky130_fd_pr__pfet_01v8_lvt_4QC8GG_1 VIN- VIN- m1_7222_1296# a_3872_2262# VSS sky130_fd_pr__pfet_01v8_lvt_4QC8GG
Xsky130_fd_pr__pfet_01v8_lvt_4QC8GG_2 VOUT VIN- m1_7222_1296# VINp VSS sky130_fd_pr__pfet_01v8_lvt_4QC8GG
Xsky130_fd_pr__nfet_01v8_lvt_8K7EBA_0 VSS m1_6338_1372# m1_7222_1296# VINp sky130_fd_pr__nfet_01v8_lvt_8K7EBA
Xsky130_fd_pr__nfet_01v8_lvt_8K7EBA_1 VSS m1_6338_1372# VSS VIN- sky130_fd_pr__nfet_01v8_lvt_8K7EBA
Xsky130_fd_pr__nfet_01v8_lvt_8K7EBA_2 VSS m1_10602_1432# VOUT VINp sky130_fd_pr__nfet_01v8_lvt_8K7EBA
Xsky130_fd_pr__nfet_01v8_lvt_8K7EBA_3 VSS a_3872_2262# m1_6338_1372# VIN- sky130_fd_pr__nfet_01v8_lvt_8K7EBA
Xsky130_fd_pr__nfet_01v8_lvt_8K7EBA_4 VSS m1_10602_1432# VSS VIN- sky130_fd_pr__nfet_01v8_lvt_8K7EBA
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_ZP6U3S c1_3269_n47100# c1_41183_n47100# m3_22126_n47200#
+ m3_n15788_n47200# m3_n34745_n47200# m3_n47383_n47200# m3_9488_n47200# c1_22226_n47100#
+ c1_n22007_n47100# c1_n40964_n47100# m3_n28426_n47200# m3_34764_n47200# c1_n9369_n47100#
+ c1_9588_n47100# m3_n41064_n47200# c1_n3050_n47100# m3_3169_n47200# c1_34864_n47100#
+ c1_n15688_n47100# c1_n34645_n47100# c1_n47283_n47100# m3_28445_n47200# m3_15807_n47200#
+ m3_n9469_n47200# m3_41083_n47200# m3_n22107_n47200# c1_28545_n47100# c1_15907_n47100#
+ c1_n28326_n47100# m3_n3150_n47200# VSUBS
X0 c1_n47283_n47100# m3_n47383_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X1 c1_41183_n47100# m3_41083_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X2 c1_n40964_n47100# m3_n41064_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X3 c1_41183_n47100# m3_41083_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X4 c1_28545_n47100# m3_28445_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X5 c1_n22007_n47100# m3_n22107_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X6 c1_34864_n47100# m3_34764_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X7 c1_n40964_n47100# m3_n41064_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X8 c1_n47283_n47100# m3_n47383_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X9 c1_34864_n47100# m3_34764_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X10 c1_n15688_n47100# m3_n15788_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X11 c1_n34645_n47100# m3_n34745_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X12 c1_15907_n47100# m3_15807_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X13 c1_n15688_n47100# m3_n15788_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X14 c1_n40964_n47100# m3_n41064_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X15 c1_9588_n47100# m3_9488_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X16 c1_n34645_n47100# m3_n34745_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X17 c1_15907_n47100# m3_15807_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X18 c1_34864_n47100# m3_34764_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X19 c1_n3050_n47100# m3_n3150_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X20 c1_n47283_n47100# m3_n47383_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X21 c1_22226_n47100# m3_22126_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X22 c1_41183_n47100# m3_41083_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X23 c1_9588_n47100# m3_9488_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X24 c1_n34645_n47100# m3_n34745_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X25 c1_n15688_n47100# m3_n15788_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X26 c1_28545_n47100# m3_28445_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X27 c1_n34645_n47100# m3_n34745_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X28 c1_15907_n47100# m3_15807_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X29 c1_28545_n47100# m3_28445_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X30 c1_15907_n47100# m3_15807_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X31 c1_n40964_n47100# m3_n41064_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X32 c1_n47283_n47100# m3_n47383_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X33 c1_15907_n47100# m3_15807_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X34 c1_3269_n47100# m3_3169_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X35 c1_n3050_n47100# m3_n3150_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X36 c1_9588_n47100# m3_9488_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X37 c1_n9369_n47100# m3_n9469_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X38 c1_28545_n47100# m3_28445_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X39 c1_41183_n47100# m3_41083_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X40 c1_n47283_n47100# m3_n47383_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X41 c1_n47283_n47100# m3_n47383_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X42 c1_15907_n47100# m3_15807_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X43 c1_9588_n47100# m3_9488_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X44 c1_n47283_n47100# m3_n47383_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X45 c1_15907_n47100# m3_15807_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X46 c1_9588_n47100# m3_9488_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X47 c1_n34645_n47100# m3_n34745_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X48 c1_n22007_n47100# m3_n22107_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X49 c1_28545_n47100# m3_28445_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X50 c1_15907_n47100# m3_15807_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X51 c1_9588_n47100# m3_9488_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X52 c1_9588_n47100# m3_9488_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X53 c1_n47283_n47100# m3_n47383_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X54 c1_28545_n47100# m3_28445_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X55 c1_n34645_n47100# m3_n34745_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X56 c1_3269_n47100# m3_3169_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X57 c1_41183_n47100# m3_41083_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X58 c1_9588_n47100# m3_9488_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X59 c1_n22007_n47100# m3_n22107_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X60 c1_n28326_n47100# m3_n28426_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X61 c1_n47283_n47100# m3_n47383_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X62 c1_28545_n47100# m3_28445_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X63 c1_n28326_n47100# m3_n28426_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X64 c1_n28326_n47100# m3_n28426_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X65 c1_22226_n47100# m3_22126_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X66 c1_n34645_n47100# m3_n34745_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X67 c1_n34645_n47100# m3_n34745_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X68 c1_n9369_n47100# m3_n9469_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X69 c1_n28326_n47100# m3_n28426_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X70 c1_15907_n47100# m3_15807_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X71 c1_3269_n47100# m3_3169_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X72 c1_n22007_n47100# m3_n22107_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X73 c1_22226_n47100# m3_22126_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X74 c1_n9369_n47100# m3_n9469_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X75 c1_9588_n47100# m3_9488_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X76 c1_n28326_n47100# m3_n28426_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X77 c1_34864_n47100# m3_34764_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X78 c1_n3050_n47100# m3_n3150_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X79 c1_22226_n47100# m3_22126_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X80 c1_3269_n47100# m3_3169_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X81 c1_n9369_n47100# m3_n9469_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X82 c1_n9369_n47100# m3_n9469_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X83 c1_41183_n47100# m3_41083_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X84 c1_22226_n47100# m3_22126_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X85 c1_n28326_n47100# m3_n28426_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X86 c1_34864_n47100# m3_34764_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X87 c1_n28326_n47100# m3_n28426_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X88 c1_34864_n47100# m3_34764_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X89 c1_n15688_n47100# m3_n15788_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X90 c1_22226_n47100# m3_22126_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X91 c1_22226_n47100# m3_22126_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X92 c1_n40964_n47100# m3_n41064_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X93 c1_n9369_n47100# m3_n9469_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X94 c1_34864_n47100# m3_34764_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X95 c1_34864_n47100# m3_34764_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X96 c1_41183_n47100# m3_41083_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X97 c1_n15688_n47100# m3_n15788_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X98 c1_n28326_n47100# m3_n28426_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X99 c1_n22007_n47100# m3_n22107_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X100 c1_n40964_n47100# m3_n41064_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X101 c1_n3050_n47100# m3_n3150_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X102 c1_n3050_n47100# m3_n3150_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X103 c1_n40964_n47100# m3_n41064_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X104 c1_3269_n47100# m3_3169_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X105 c1_n47283_n47100# m3_n47383_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X106 c1_n47283_n47100# m3_n47383_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X107 c1_15907_n47100# m3_15807_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X108 c1_28545_n47100# m3_28445_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X109 c1_n40964_n47100# m3_n41064_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X110 c1_41183_n47100# m3_41083_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X111 c1_n22007_n47100# m3_n22107_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X112 c1_n15688_n47100# m3_n15788_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X113 c1_n40964_n47100# m3_n41064_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X114 c1_28545_n47100# m3_28445_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X115 c1_3269_n47100# m3_3169_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X116 c1_9588_n47100# m3_9488_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X117 c1_n15688_n47100# m3_n15788_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X118 c1_34864_n47100# m3_34764_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X119 c1_n15688_n47100# m3_n15788_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X120 c1_n3050_n47100# m3_n3150_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X121 c1_41183_n47100# m3_41083_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X122 c1_n3050_n47100# m3_n3150_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X123 c1_n3050_n47100# m3_n3150_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X124 c1_n15688_n47100# m3_n15788_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X125 c1_9588_n47100# m3_9488_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X126 c1_n22007_n47100# m3_n22107_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X127 c1_28545_n47100# m3_28445_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X128 c1_n3050_n47100# m3_n3150_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X129 c1_n3050_n47100# m3_n3150_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X130 c1_n3050_n47100# m3_n3150_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X131 c1_22226_n47100# m3_22126_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X132 c1_n34645_n47100# m3_n34745_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X133 c1_n34645_n47100# m3_n34745_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X134 c1_28545_n47100# m3_28445_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X135 c1_28545_n47100# m3_28445_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X136 c1_15907_n47100# m3_15807_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X137 c1_n40964_n47100# m3_n41064_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X138 c1_41183_n47100# m3_41083_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X139 c1_3269_n47100# m3_3169_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X140 c1_34864_n47100# m3_34764_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X141 c1_n15688_n47100# m3_n15788_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X142 c1_9588_n47100# m3_9488_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X143 c1_n22007_n47100# m3_n22107_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X144 c1_n47283_n47100# m3_n47383_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X145 c1_15907_n47100# m3_15807_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X146 c1_n47283_n47100# m3_n47383_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X147 c1_41183_n47100# m3_41083_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X148 c1_41183_n47100# m3_41083_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X149 c1_22226_n47100# m3_22126_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X150 c1_n34645_n47100# m3_n34745_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X151 c1_n22007_n47100# m3_n22107_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X152 c1_28545_n47100# m3_28445_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X153 c1_n9369_n47100# m3_n9469_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X154 c1_n22007_n47100# m3_n22107_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X155 c1_9588_n47100# m3_9488_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X156 c1_n40964_n47100# m3_n41064_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X157 c1_n47283_n47100# m3_n47383_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X158 c1_15907_n47100# m3_15807_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X159 c1_n34645_n47100# m3_n34745_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X160 c1_n34645_n47100# m3_n34745_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X161 c1_9588_n47100# m3_9488_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X162 c1_3269_n47100# m3_3169_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X163 c1_n28326_n47100# m3_n28426_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X164 c1_22226_n47100# m3_22126_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X165 c1_n47283_n47100# m3_n47383_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X166 c1_9588_n47100# m3_9488_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X167 c1_22226_n47100# m3_22126_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X168 c1_n34645_n47100# m3_n34745_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X169 c1_41183_n47100# m3_41083_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X170 c1_n9369_n47100# m3_n9469_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X171 c1_28545_n47100# m3_28445_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X172 c1_n9369_n47100# m3_n9469_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X173 c1_3269_n47100# m3_3169_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X174 c1_34864_n47100# m3_34764_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X175 c1_n15688_n47100# m3_n15788_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X176 c1_15907_n47100# m3_15807_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X177 c1_3269_n47100# m3_3169_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X178 c1_n28326_n47100# m3_n28426_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X179 c1_41183_n47100# m3_41083_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X180 c1_n9369_n47100# m3_n9469_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X181 c1_n22007_n47100# m3_n22107_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X182 c1_22226_n47100# m3_22126_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X183 c1_n9369_n47100# m3_n9469_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X184 c1_n15688_n47100# m3_n15788_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X185 c1_n3050_n47100# m3_n3150_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X186 c1_22226_n47100# m3_22126_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X187 c1_n34645_n47100# m3_n34745_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X188 c1_n22007_n47100# m3_n22107_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X189 c1_15907_n47100# m3_15807_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X190 c1_3269_n47100# m3_3169_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X191 c1_41183_n47100# m3_41083_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X192 c1_n40964_n47100# m3_n41064_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X193 c1_n28326_n47100# m3_n28426_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X194 c1_n22007_n47100# m3_n22107_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X195 c1_n22007_n47100# m3_n22107_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X196 c1_3269_n47100# m3_3169_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X197 c1_n28326_n47100# m3_n28426_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X198 c1_22226_n47100# m3_22126_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X199 c1_n28326_n47100# m3_n28426_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X200 c1_34864_n47100# m3_34764_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X201 c1_n3050_n47100# m3_n3150_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X202 c1_n28326_n47100# m3_n28426_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X203 c1_n15688_n47100# m3_n15788_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X204 c1_n15688_n47100# m3_n15788_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X205 c1_n40964_n47100# m3_n41064_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X206 c1_n9369_n47100# m3_n9469_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X207 c1_34864_n47100# m3_34764_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X208 c1_n3050_n47100# m3_n3150_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X209 c1_n22007_n47100# m3_n22107_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X210 c1_22226_n47100# m3_22126_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X211 c1_n40964_n47100# m3_n41064_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X212 c1_3269_n47100# m3_3169_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X213 c1_28545_n47100# m3_28445_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X214 c1_n9369_n47100# m3_n9469_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X215 c1_n28326_n47100# m3_n28426_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X216 c1_34864_n47100# m3_34764_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X217 c1_n40964_n47100# m3_n41064_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X218 c1_34864_n47100# m3_34764_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X219 c1_n15688_n47100# m3_n15788_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X220 c1_n3050_n47100# m3_n3150_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X221 c1_3269_n47100# m3_3169_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X222 c1_n9369_n47100# m3_n9469_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X223 c1_3269_n47100# m3_3169_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X224 c1_n9369_n47100# m3_n9469_n47200# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
.ends

.subckt cap225_layout VIN VOUT VSUBS
Xsky130_fd_pr__cap_mim_m3_1_ZP6U3S_0 VIN VIN VOUT VOUT VOUT VOUT VOUT VIN VIN VIN
+ VOUT VOUT VIN VIN VOUT VIN VOUT VIN VIN VIN VIN VOUT VOUT VOUT VOUT VOUT VIN VIN
+ VIN VOUT VSUBS sky130_fd_pr__cap_mim_m3_1_ZP6U3S
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_4QDPGG w_n231_n8219# a_n35_n8097# a_35_n8000#
+ a_n93_n8000# VSUBS
X0 a_35_n8000# a_n35_n8097# a_n93_n8000# w_n231_n8219# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+07u l=350000u
.ends

.subckt pmos20 G D B S VSUBS
Xsky130_fd_pr__pfet_01v8_lvt_4QDPGG_0[0] B G S D sky130_fd_pr__pfet_01v8_lvt_4QDPGG_0[0]/VSUBS
+ sky130_fd_pr__pfet_01v8_lvt_4QDPGG
Xsky130_fd_pr__pfet_01v8_lvt_4QDPGG_0[1] B G S D sky130_fd_pr__pfet_01v8_lvt_4QDPGG_0[1]/VSUBS
+ sky130_fd_pr__pfet_01v8_lvt_4QDPGG
Xsky130_fd_pr__pfet_01v8_lvt_4QDPGG_0[2] B G S D sky130_fd_pr__pfet_01v8_lvt_4QDPGG_0[2]/VSUBS
+ sky130_fd_pr__pfet_01v8_lvt_4QDPGG
Xsky130_fd_pr__pfet_01v8_lvt_4QDPGG_0[3] B G S D sky130_fd_pr__pfet_01v8_lvt_4QDPGG_0[3]/VSUBS
+ sky130_fd_pr__pfet_01v8_lvt_4QDPGG
Xsky130_fd_pr__pfet_01v8_lvt_4QDPGG_0[4] B G S D sky130_fd_pr__pfet_01v8_lvt_4QDPGG_0[4]/VSUBS
+ sky130_fd_pr__pfet_01v8_lvt_4QDPGG
Xsky130_fd_pr__pfet_01v8_lvt_4QDPGG_0[5] B G S D sky130_fd_pr__pfet_01v8_lvt_4QDPGG_0[5]/VSUBS
+ sky130_fd_pr__pfet_01v8_lvt_4QDPGG
Xsky130_fd_pr__pfet_01v8_lvt_4QDPGG_0[6] B G S D sky130_fd_pr__pfet_01v8_lvt_4QDPGG_0[6]/VSUBS
+ sky130_fd_pr__pfet_01v8_lvt_4QDPGG
Xsky130_fd_pr__pfet_01v8_lvt_4QDPGG_0[7] B G S D sky130_fd_pr__pfet_01v8_lvt_4QDPGG_0[7]/VSUBS
+ sky130_fd_pr__pfet_01v8_lvt_4QDPGG
Xsky130_fd_pr__pfet_01v8_lvt_4QDPGG_0[8] B G S D sky130_fd_pr__pfet_01v8_lvt_4QDPGG_0[8]/VSUBS
+ sky130_fd_pr__pfet_01v8_lvt_4QDPGG
Xsky130_fd_pr__pfet_01v8_lvt_4QDPGG_0[9] B G S D sky130_fd_pr__pfet_01v8_lvt_4QDPGG_0[9]/VSUBS
+ sky130_fd_pr__pfet_01v8_lvt_4QDPGG
Xsky130_fd_pr__pfet_01v8_lvt_4QDPGG_0[10] B G S D sky130_fd_pr__pfet_01v8_lvt_4QDPGG_0[10]/VSUBS
+ sky130_fd_pr__pfet_01v8_lvt_4QDPGG
Xsky130_fd_pr__pfet_01v8_lvt_4QDPGG_0[11] B G S D sky130_fd_pr__pfet_01v8_lvt_4QDPGG_0[11]/VSUBS
+ sky130_fd_pr__pfet_01v8_lvt_4QDPGG
Xsky130_fd_pr__pfet_01v8_lvt_4QDPGG_0[12] B G S D sky130_fd_pr__pfet_01v8_lvt_4QDPGG_0[12]/VSUBS
+ sky130_fd_pr__pfet_01v8_lvt_4QDPGG
Xsky130_fd_pr__pfet_01v8_lvt_4QDPGG_0[13] B G S D sky130_fd_pr__pfet_01v8_lvt_4QDPGG_0[13]/VSUBS
+ sky130_fd_pr__pfet_01v8_lvt_4QDPGG
Xsky130_fd_pr__pfet_01v8_lvt_4QDPGG_0[14] B G S D sky130_fd_pr__pfet_01v8_lvt_4QDPGG_0[14]/VSUBS
+ sky130_fd_pr__pfet_01v8_lvt_4QDPGG
Xsky130_fd_pr__pfet_01v8_lvt_4QDPGG_0[15] B G S D sky130_fd_pr__pfet_01v8_lvt_4QDPGG_0[15]/VSUBS
+ sky130_fd_pr__pfet_01v8_lvt_4QDPGG
Xsky130_fd_pr__pfet_01v8_lvt_4QDPGG_0[16] B G S D sky130_fd_pr__pfet_01v8_lvt_4QDPGG_0[16]/VSUBS
+ sky130_fd_pr__pfet_01v8_lvt_4QDPGG
Xsky130_fd_pr__pfet_01v8_lvt_4QDPGG_0[17] B G S D sky130_fd_pr__pfet_01v8_lvt_4QDPGG_0[17]/VSUBS
+ sky130_fd_pr__pfet_01v8_lvt_4QDPGG
Xsky130_fd_pr__pfet_01v8_lvt_4QDPGG_0[18] B G S D VSUBS sky130_fd_pr__pfet_01v8_lvt_4QDPGG
Xsky130_fd_pr__pfet_01v8_lvt_4QDPGG_0[19] B G S D sky130_fd_pr__pfet_01v8_lvt_4QDPGG_0[19]/VSUBS
+ sky130_fd_pr__pfet_01v8_lvt_4QDPGG
.ends

.subckt pmos40 pmos20_0[1]/S pmos20_0[1]/G pmos20_0[1]/B pmos20_0[1]/D VSUBS
Xpmos20_0[0] pmos20_0[1]/G pmos20_0[1]/D pmos20_0[1]/B pmos20_0[1]/S VSUBS pmos20
Xpmos20_0[1] pmos20_0[1]/G pmos20_0[1]/D pmos20_0[1]/B pmos20_0[1]/S pmos20_0[1]/VSUBS
+ pmos20
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_BPY4AF a_35_n8000# a_n35_n8088# w_n231_n8210#
+ a_n93_n8000#
X0 a_35_n8000# a_n35_n8088# a_n93_n8000# w_n231_n8210# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+07u l=350000u
.ends

.subckt nmos20 G B D S
Xsky130_fd_pr__nfet_01v8_lvt_BPY4AF_0[0] S G B D sky130_fd_pr__nfet_01v8_lvt_BPY4AF
Xsky130_fd_pr__nfet_01v8_lvt_BPY4AF_0[1] S G B D sky130_fd_pr__nfet_01v8_lvt_BPY4AF
Xsky130_fd_pr__nfet_01v8_lvt_BPY4AF_0[2] S G B D sky130_fd_pr__nfet_01v8_lvt_BPY4AF
Xsky130_fd_pr__nfet_01v8_lvt_BPY4AF_0[3] S G B D sky130_fd_pr__nfet_01v8_lvt_BPY4AF
Xsky130_fd_pr__nfet_01v8_lvt_BPY4AF_0[4] S G B D sky130_fd_pr__nfet_01v8_lvt_BPY4AF
Xsky130_fd_pr__nfet_01v8_lvt_BPY4AF_0[5] S G B D sky130_fd_pr__nfet_01v8_lvt_BPY4AF
Xsky130_fd_pr__nfet_01v8_lvt_BPY4AF_0[6] S G B D sky130_fd_pr__nfet_01v8_lvt_BPY4AF
Xsky130_fd_pr__nfet_01v8_lvt_BPY4AF_0[7] S G B D sky130_fd_pr__nfet_01v8_lvt_BPY4AF
Xsky130_fd_pr__nfet_01v8_lvt_BPY4AF_0[8] S G B D sky130_fd_pr__nfet_01v8_lvt_BPY4AF
Xsky130_fd_pr__nfet_01v8_lvt_BPY4AF_0[9] S G B D sky130_fd_pr__nfet_01v8_lvt_BPY4AF
Xsky130_fd_pr__nfet_01v8_lvt_BPY4AF_0[10] S G B D sky130_fd_pr__nfet_01v8_lvt_BPY4AF
Xsky130_fd_pr__nfet_01v8_lvt_BPY4AF_0[11] S G B D sky130_fd_pr__nfet_01v8_lvt_BPY4AF
Xsky130_fd_pr__nfet_01v8_lvt_BPY4AF_0[12] S G B D sky130_fd_pr__nfet_01v8_lvt_BPY4AF
Xsky130_fd_pr__nfet_01v8_lvt_BPY4AF_0[13] S G B D sky130_fd_pr__nfet_01v8_lvt_BPY4AF
Xsky130_fd_pr__nfet_01v8_lvt_BPY4AF_0[14] S G B D sky130_fd_pr__nfet_01v8_lvt_BPY4AF
Xsky130_fd_pr__nfet_01v8_lvt_BPY4AF_0[15] S G B D sky130_fd_pr__nfet_01v8_lvt_BPY4AF
Xsky130_fd_pr__nfet_01v8_lvt_BPY4AF_0[16] S G B D sky130_fd_pr__nfet_01v8_lvt_BPY4AF
Xsky130_fd_pr__nfet_01v8_lvt_BPY4AF_0[17] S G B D sky130_fd_pr__nfet_01v8_lvt_BPY4AF
Xsky130_fd_pr__nfet_01v8_lvt_BPY4AF_0[18] S G B D sky130_fd_pr__nfet_01v8_lvt_BPY4AF
Xsky130_fd_pr__nfet_01v8_lvt_BPY4AF_0[19] S G B D sky130_fd_pr__nfet_01v8_lvt_BPY4AF
.ends

.subckt recitifer_layout VINN VIN1 VINP VSS
Xpmos20_0 VINN VIN1 VINP VINP VSS pmos20
Xpmos20_1 VINP VIN1 VINN VINN VSS pmos20
Xnmos20_0 VINN VSS VINP VSS nmos20
Xnmos20_1 VINP VSS VINN VSS nmos20
.ends

.subckt RX_layout VIN2 VIN1 recitifer_layout_0/VINP VOUT_C recitifer_layout_0/VINN
+ VSS
Xcap225_layout_0 VIN2 VSS VSS cap225_layout
Xpmos40_0 VIN1 VOUT_C VIN2 VIN2 VSS pmos40
Xrecitifer_layout_0 recitifer_layout_0/VINN VIN1 recitifer_layout_0/VINP VSS recitifer_layout
Xpmos40_1 VIN2 VOUT_C VIN2 pmos40_1/pmos20_0[1]/D VSS pmos40
.ends

.subckt FINAL RX_layout_0/recitifer_layout_0/VINP RX_layout_0/recitifer_layout_0/VINN
+ VSUBS
XComparator_jafar_0 VSUBS RX_layout_0/VIN1 RX_layout_0/VIN2 RX_layout_0/VOUT_C Comparator_jafar
XRX_layout_0 RX_layout_0/VIN2 RX_layout_0/VIN1 RX_layout_0/recitifer_layout_0/VINP
+ RX_layout_0/VOUT_C RX_layout_0/recitifer_layout_0/VINN VSUBS RX_layout
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_NBPZFR m3_n24306_n24190# m3_6089_n24190# m3_n12148_n24190#
+ m3_10_n24190# c1_6189_n24090# m3_n6069_n24190# c1_n5969_n24090# c1_n18127_n24090#
+ c1_n24206_n24090# c1_n12048_n24090# m3_18247_n24190# m3_12168_n24190# c1_18347_n24090#
+ c1_12268_n24090# c1_110_n24090# m3_n18227_n24190# VSUBS
X0 c1_12268_n24090# m3_12168_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X1 c1_n5969_n24090# m3_n6069_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X2 c1_6189_n24090# m3_6089_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X3 c1_110_n24090# m3_10_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X4 c1_n24206_n24090# m3_n24306_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X5 c1_n24206_n24090# m3_n24306_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X6 c1_n18127_n24090# m3_n18227_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X7 c1_110_n24090# m3_10_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X8 c1_12268_n24090# m3_12168_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X9 c1_n24206_n24090# m3_n24306_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X10 c1_n5969_n24090# m3_n6069_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X11 c1_n18127_n24090# m3_n18227_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X12 c1_6189_n24090# m3_6089_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X13 c1_n12048_n24090# m3_n12148_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X14 c1_12268_n24090# m3_12168_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X15 c1_110_n24090# m3_10_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X16 c1_18347_n24090# m3_18247_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X17 c1_12268_n24090# m3_12168_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X18 c1_110_n24090# m3_10_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X19 c1_n24206_n24090# m3_n24306_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X20 c1_110_n24090# m3_10_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X21 c1_18347_n24090# m3_18247_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X22 c1_n24206_n24090# m3_n24306_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X23 c1_6189_n24090# m3_6089_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X24 c1_12268_n24090# m3_12168_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X25 c1_n24206_n24090# m3_n24306_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X26 c1_n12048_n24090# m3_n12148_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X27 c1_12268_n24090# m3_12168_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X28 c1_n24206_n24090# m3_n24306_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X29 c1_n18127_n24090# m3_n18227_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X30 c1_n18127_n24090# m3_n18227_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X31 c1_n12048_n24090# m3_n12148_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X32 c1_110_n24090# m3_10_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X33 c1_18347_n24090# m3_18247_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X34 c1_110_n24090# m3_10_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X35 c1_18347_n24090# m3_18247_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X36 c1_n12048_n24090# m3_n12148_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X37 c1_6189_n24090# m3_6089_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X38 c1_6189_n24090# m3_6089_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X39 c1_6189_n24090# m3_6089_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X40 c1_6189_n24090# m3_6089_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X41 c1_n5969_n24090# m3_n6069_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X42 c1_n18127_n24090# m3_n18227_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X43 c1_110_n24090# m3_10_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X44 c1_18347_n24090# m3_18247_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X45 c1_n24206_n24090# m3_n24306_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X46 c1_n12048_n24090# m3_n12148_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X47 c1_n5969_n24090# m3_n6069_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X48 c1_n12048_n24090# m3_n12148_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X49 c1_n12048_n24090# m3_n12148_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X50 c1_12268_n24090# m3_12168_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X51 c1_n5969_n24090# m3_n6069_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X52 c1_n5969_n24090# m3_n6069_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X53 c1_n18127_n24090# m3_n18227_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X54 c1_6189_n24090# m3_6089_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X55 c1_n5969_n24090# m3_n6069_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X56 c1_n18127_n24090# m3_n18227_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X57 c1_n12048_n24090# m3_n12148_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X58 c1_18347_n24090# m3_18247_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X59 c1_12268_n24090# m3_12168_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X60 c1_n18127_n24090# m3_n18227_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X61 c1_18347_n24090# m3_18247_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X62 c1_n5969_n24090# m3_n6069_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
X63 c1_18347_n24090# m3_18247_n24190# sky130_fd_pr__cap_mim_m3_1 l=2.88e+07u w=2.88e+07u
.ends

.subckt cap107_layout VIN VOUT VSUBS
Xsky130_fd_pr__cap_mim_m3_1_NBPZFR_0 VOUT VOUT VOUT VOUT VIN VOUT VIN VIN VIN VIN
+ VOUT VOUT VIN VIN VIN VOUT VSUBS sky130_fd_pr__cap_mim_m3_1_NBPZFR
.ends


* Top level circuit FINAL_without_ind

XFINAL_0 VINP VINN VSUBS FINAL
Xcap107_layout_0 VINP VINN VSUBS cap107_layout
.end

