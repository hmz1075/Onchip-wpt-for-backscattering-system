magic
tech sky130A
magscale 1 2
timestamp 1634724870
<< error_p >>
rect -39194 15050 -39134 20950
rect -39114 15050 -39054 20950
rect -33175 15050 -33115 20950
rect -33095 15050 -33035 20950
rect -27156 15050 -27096 20950
rect -27076 15050 -27016 20950
rect -21137 15050 -21077 20950
rect -21057 15050 -20997 20950
rect -15118 15050 -15058 20950
rect -15038 15050 -14978 20950
rect -9099 15050 -9039 20950
rect -9019 15050 -8959 20950
rect -3080 15050 -3020 20950
rect -3000 15050 -2940 20950
rect 2939 15050 2999 20950
rect 3019 15050 3079 20950
rect 8958 15050 9018 20950
rect 9038 15050 9098 20950
rect 14977 15050 15037 20950
rect 15057 15050 15117 20950
rect 20996 15050 21056 20950
rect 21076 15050 21136 20950
rect 27015 15050 27075 20950
rect 27095 15050 27155 20950
rect 33034 15050 33094 20950
rect 33114 15050 33174 20950
rect 39053 15050 39113 20950
rect 39133 15050 39193 20950
rect -39194 9050 -39134 14950
rect -39114 9050 -39054 14950
rect -33175 9050 -33115 14950
rect -33095 9050 -33035 14950
rect -27156 9050 -27096 14950
rect -27076 9050 -27016 14950
rect -21137 9050 -21077 14950
rect -21057 9050 -20997 14950
rect -15118 9050 -15058 14950
rect -15038 9050 -14978 14950
rect -9099 9050 -9039 14950
rect -9019 9050 -8959 14950
rect -3080 9050 -3020 14950
rect -3000 9050 -2940 14950
rect 2939 9050 2999 14950
rect 3019 9050 3079 14950
rect 8958 9050 9018 14950
rect 9038 9050 9098 14950
rect 14977 9050 15037 14950
rect 15057 9050 15117 14950
rect 20996 9050 21056 14950
rect 21076 9050 21136 14950
rect 27015 9050 27075 14950
rect 27095 9050 27155 14950
rect 33034 9050 33094 14950
rect 33114 9050 33174 14950
rect 39053 9050 39113 14950
rect 39133 9050 39193 14950
rect -39194 3050 -39134 8950
rect -39114 3050 -39054 8950
rect -33175 3050 -33115 8950
rect -33095 3050 -33035 8950
rect -27156 3050 -27096 8950
rect -27076 3050 -27016 8950
rect -21137 3050 -21077 8950
rect -21057 3050 -20997 8950
rect -15118 3050 -15058 8950
rect -15038 3050 -14978 8950
rect -9099 3050 -9039 8950
rect -9019 3050 -8959 8950
rect -3080 3050 -3020 8950
rect -3000 3050 -2940 8950
rect 2939 3050 2999 8950
rect 3019 3050 3079 8950
rect 8958 3050 9018 8950
rect 9038 3050 9098 8950
rect 14977 3050 15037 8950
rect 15057 3050 15117 8950
rect 20996 3050 21056 8950
rect 21076 3050 21136 8950
rect 27015 3050 27075 8950
rect 27095 3050 27155 8950
rect 33034 3050 33094 8950
rect 33114 3050 33174 8950
rect 39053 3050 39113 8950
rect 39133 3050 39193 8950
rect -39194 -2950 -39134 2950
rect -39114 -2950 -39054 2950
rect -33175 -2950 -33115 2950
rect -33095 -2950 -33035 2950
rect -27156 -2950 -27096 2950
rect -27076 -2950 -27016 2950
rect -21137 -2950 -21077 2950
rect -21057 -2950 -20997 2950
rect -15118 -2950 -15058 2950
rect -15038 -2950 -14978 2950
rect -9099 -2950 -9039 2950
rect -9019 -2950 -8959 2950
rect -3080 -2950 -3020 2950
rect -3000 -2950 -2940 2950
rect 2939 -2950 2999 2950
rect 3019 -2950 3079 2950
rect 8958 -2950 9018 2950
rect 9038 -2950 9098 2950
rect 14977 -2950 15037 2950
rect 15057 -2950 15117 2950
rect 20996 -2950 21056 2950
rect 21076 -2950 21136 2950
rect 27015 -2950 27075 2950
rect 27095 -2950 27155 2950
rect 33034 -2950 33094 2950
rect 33114 -2950 33174 2950
rect 39053 -2950 39113 2950
rect 39133 -2950 39193 2950
rect -39194 -8950 -39134 -3050
rect -39114 -8950 -39054 -3050
rect -33175 -8950 -33115 -3050
rect -33095 -8950 -33035 -3050
rect -27156 -8950 -27096 -3050
rect -27076 -8950 -27016 -3050
rect -21137 -8950 -21077 -3050
rect -21057 -8950 -20997 -3050
rect -15118 -8950 -15058 -3050
rect -15038 -8950 -14978 -3050
rect -9099 -8950 -9039 -3050
rect -9019 -8950 -8959 -3050
rect -3080 -8950 -3020 -3050
rect -3000 -8950 -2940 -3050
rect 2939 -8950 2999 -3050
rect 3019 -8950 3079 -3050
rect 8958 -8950 9018 -3050
rect 9038 -8950 9098 -3050
rect 14977 -8950 15037 -3050
rect 15057 -8950 15117 -3050
rect 20996 -8950 21056 -3050
rect 21076 -8950 21136 -3050
rect 27015 -8950 27075 -3050
rect 27095 -8950 27155 -3050
rect 33034 -8950 33094 -3050
rect 33114 -8950 33174 -3050
rect 39053 -8950 39113 -3050
rect 39133 -8950 39193 -3050
rect -39194 -14950 -39134 -9050
rect -39114 -14950 -39054 -9050
rect -33175 -14950 -33115 -9050
rect -33095 -14950 -33035 -9050
rect -27156 -14950 -27096 -9050
rect -27076 -14950 -27016 -9050
rect -21137 -14950 -21077 -9050
rect -21057 -14950 -20997 -9050
rect -15118 -14950 -15058 -9050
rect -15038 -14950 -14978 -9050
rect -9099 -14950 -9039 -9050
rect -9019 -14950 -8959 -9050
rect -3080 -14950 -3020 -9050
rect -3000 -14950 -2940 -9050
rect 2939 -14950 2999 -9050
rect 3019 -14950 3079 -9050
rect 8958 -14950 9018 -9050
rect 9038 -14950 9098 -9050
rect 14977 -14950 15037 -9050
rect 15057 -14950 15117 -9050
rect 20996 -14950 21056 -9050
rect 21076 -14950 21136 -9050
rect 27015 -14950 27075 -9050
rect 27095 -14950 27155 -9050
rect 33034 -14950 33094 -9050
rect 33114 -14950 33174 -9050
rect 39053 -14950 39113 -9050
rect 39133 -14950 39193 -9050
rect -39194 -20950 -39134 -15050
rect -39114 -20950 -39054 -15050
rect -33175 -20950 -33115 -15050
rect -33095 -20950 -33035 -15050
rect -27156 -20950 -27096 -15050
rect -27076 -20950 -27016 -15050
rect -21137 -20950 -21077 -15050
rect -21057 -20950 -20997 -15050
rect -15118 -20950 -15058 -15050
rect -15038 -20950 -14978 -15050
rect -9099 -20950 -9039 -15050
rect -9019 -20950 -8959 -15050
rect -3080 -20950 -3020 -15050
rect -3000 -20950 -2940 -15050
rect 2939 -20950 2999 -15050
rect 3019 -20950 3079 -15050
rect 8958 -20950 9018 -15050
rect 9038 -20950 9098 -15050
rect 14977 -20950 15037 -15050
rect 15057 -20950 15117 -15050
rect 20996 -20950 21056 -15050
rect 21076 -20950 21136 -15050
rect 27015 -20950 27075 -15050
rect 27095 -20950 27155 -15050
rect 33034 -20950 33094 -15050
rect 33114 -20950 33174 -15050
rect 39053 -20950 39113 -15050
rect 39133 -20950 39193 -15050
<< metal3 >>
rect -45133 20922 -39134 20950
rect -45133 15078 -39218 20922
rect -39154 15078 -39134 20922
rect -45133 15050 -39134 15078
rect -39114 20922 -33115 20950
rect -39114 15078 -33199 20922
rect -33135 15078 -33115 20922
rect -39114 15050 -33115 15078
rect -33095 20922 -27096 20950
rect -33095 15078 -27180 20922
rect -27116 15078 -27096 20922
rect -33095 15050 -27096 15078
rect -27076 20922 -21077 20950
rect -27076 15078 -21161 20922
rect -21097 15078 -21077 20922
rect -27076 15050 -21077 15078
rect -21057 20922 -15058 20950
rect -21057 15078 -15142 20922
rect -15078 15078 -15058 20922
rect -21057 15050 -15058 15078
rect -15038 20922 -9039 20950
rect -15038 15078 -9123 20922
rect -9059 15078 -9039 20922
rect -15038 15050 -9039 15078
rect -9019 20922 -3020 20950
rect -9019 15078 -3104 20922
rect -3040 15078 -3020 20922
rect -9019 15050 -3020 15078
rect -3000 20922 2999 20950
rect -3000 15078 2915 20922
rect 2979 15078 2999 20922
rect -3000 15050 2999 15078
rect 3019 20922 9018 20950
rect 3019 15078 8934 20922
rect 8998 15078 9018 20922
rect 3019 15050 9018 15078
rect 9038 20922 15037 20950
rect 9038 15078 14953 20922
rect 15017 15078 15037 20922
rect 9038 15050 15037 15078
rect 15057 20922 21056 20950
rect 15057 15078 20972 20922
rect 21036 15078 21056 20922
rect 15057 15050 21056 15078
rect 21076 20922 27075 20950
rect 21076 15078 26991 20922
rect 27055 15078 27075 20922
rect 21076 15050 27075 15078
rect 27095 20922 33094 20950
rect 27095 15078 33010 20922
rect 33074 15078 33094 20922
rect 27095 15050 33094 15078
rect 33114 20922 39113 20950
rect 33114 15078 39029 20922
rect 39093 15078 39113 20922
rect 33114 15050 39113 15078
rect 39133 20922 45132 20950
rect 39133 15078 45048 20922
rect 45112 15078 45132 20922
rect 39133 15050 45132 15078
rect -45133 14922 -39134 14950
rect -45133 9078 -39218 14922
rect -39154 9078 -39134 14922
rect -45133 9050 -39134 9078
rect -39114 14922 -33115 14950
rect -39114 9078 -33199 14922
rect -33135 9078 -33115 14922
rect -39114 9050 -33115 9078
rect -33095 14922 -27096 14950
rect -33095 9078 -27180 14922
rect -27116 9078 -27096 14922
rect -33095 9050 -27096 9078
rect -27076 14922 -21077 14950
rect -27076 9078 -21161 14922
rect -21097 9078 -21077 14922
rect -27076 9050 -21077 9078
rect -21057 14922 -15058 14950
rect -21057 9078 -15142 14922
rect -15078 9078 -15058 14922
rect -21057 9050 -15058 9078
rect -15038 14922 -9039 14950
rect -15038 9078 -9123 14922
rect -9059 9078 -9039 14922
rect -15038 9050 -9039 9078
rect -9019 14922 -3020 14950
rect -9019 9078 -3104 14922
rect -3040 9078 -3020 14922
rect -9019 9050 -3020 9078
rect -3000 14922 2999 14950
rect -3000 9078 2915 14922
rect 2979 9078 2999 14922
rect -3000 9050 2999 9078
rect 3019 14922 9018 14950
rect 3019 9078 8934 14922
rect 8998 9078 9018 14922
rect 3019 9050 9018 9078
rect 9038 14922 15037 14950
rect 9038 9078 14953 14922
rect 15017 9078 15037 14922
rect 9038 9050 15037 9078
rect 15057 14922 21056 14950
rect 15057 9078 20972 14922
rect 21036 9078 21056 14922
rect 15057 9050 21056 9078
rect 21076 14922 27075 14950
rect 21076 9078 26991 14922
rect 27055 9078 27075 14922
rect 21076 9050 27075 9078
rect 27095 14922 33094 14950
rect 27095 9078 33010 14922
rect 33074 9078 33094 14922
rect 27095 9050 33094 9078
rect 33114 14922 39113 14950
rect 33114 9078 39029 14922
rect 39093 9078 39113 14922
rect 33114 9050 39113 9078
rect 39133 14922 45132 14950
rect 39133 9078 45048 14922
rect 45112 9078 45132 14922
rect 39133 9050 45132 9078
rect -45133 8922 -39134 8950
rect -45133 3078 -39218 8922
rect -39154 3078 -39134 8922
rect -45133 3050 -39134 3078
rect -39114 8922 -33115 8950
rect -39114 3078 -33199 8922
rect -33135 3078 -33115 8922
rect -39114 3050 -33115 3078
rect -33095 8922 -27096 8950
rect -33095 3078 -27180 8922
rect -27116 3078 -27096 8922
rect -33095 3050 -27096 3078
rect -27076 8922 -21077 8950
rect -27076 3078 -21161 8922
rect -21097 3078 -21077 8922
rect -27076 3050 -21077 3078
rect -21057 8922 -15058 8950
rect -21057 3078 -15142 8922
rect -15078 3078 -15058 8922
rect -21057 3050 -15058 3078
rect -15038 8922 -9039 8950
rect -15038 3078 -9123 8922
rect -9059 3078 -9039 8922
rect -15038 3050 -9039 3078
rect -9019 8922 -3020 8950
rect -9019 3078 -3104 8922
rect -3040 3078 -3020 8922
rect -9019 3050 -3020 3078
rect -3000 8922 2999 8950
rect -3000 3078 2915 8922
rect 2979 3078 2999 8922
rect -3000 3050 2999 3078
rect 3019 8922 9018 8950
rect 3019 3078 8934 8922
rect 8998 3078 9018 8922
rect 3019 3050 9018 3078
rect 9038 8922 15037 8950
rect 9038 3078 14953 8922
rect 15017 3078 15037 8922
rect 9038 3050 15037 3078
rect 15057 8922 21056 8950
rect 15057 3078 20972 8922
rect 21036 3078 21056 8922
rect 15057 3050 21056 3078
rect 21076 8922 27075 8950
rect 21076 3078 26991 8922
rect 27055 3078 27075 8922
rect 21076 3050 27075 3078
rect 27095 8922 33094 8950
rect 27095 3078 33010 8922
rect 33074 3078 33094 8922
rect 27095 3050 33094 3078
rect 33114 8922 39113 8950
rect 33114 3078 39029 8922
rect 39093 3078 39113 8922
rect 33114 3050 39113 3078
rect 39133 8922 45132 8950
rect 39133 3078 45048 8922
rect 45112 3078 45132 8922
rect 39133 3050 45132 3078
rect -45133 2922 -39134 2950
rect -45133 -2922 -39218 2922
rect -39154 -2922 -39134 2922
rect -45133 -2950 -39134 -2922
rect -39114 2922 -33115 2950
rect -39114 -2922 -33199 2922
rect -33135 -2922 -33115 2922
rect -39114 -2950 -33115 -2922
rect -33095 2922 -27096 2950
rect -33095 -2922 -27180 2922
rect -27116 -2922 -27096 2922
rect -33095 -2950 -27096 -2922
rect -27076 2922 -21077 2950
rect -27076 -2922 -21161 2922
rect -21097 -2922 -21077 2922
rect -27076 -2950 -21077 -2922
rect -21057 2922 -15058 2950
rect -21057 -2922 -15142 2922
rect -15078 -2922 -15058 2922
rect -21057 -2950 -15058 -2922
rect -15038 2922 -9039 2950
rect -15038 -2922 -9123 2922
rect -9059 -2922 -9039 2922
rect -15038 -2950 -9039 -2922
rect -9019 2922 -3020 2950
rect -9019 -2922 -3104 2922
rect -3040 -2922 -3020 2922
rect -9019 -2950 -3020 -2922
rect -3000 2922 2999 2950
rect -3000 -2922 2915 2922
rect 2979 -2922 2999 2922
rect -3000 -2950 2999 -2922
rect 3019 2922 9018 2950
rect 3019 -2922 8934 2922
rect 8998 -2922 9018 2922
rect 3019 -2950 9018 -2922
rect 9038 2922 15037 2950
rect 9038 -2922 14953 2922
rect 15017 -2922 15037 2922
rect 9038 -2950 15037 -2922
rect 15057 2922 21056 2950
rect 15057 -2922 20972 2922
rect 21036 -2922 21056 2922
rect 15057 -2950 21056 -2922
rect 21076 2922 27075 2950
rect 21076 -2922 26991 2922
rect 27055 -2922 27075 2922
rect 21076 -2950 27075 -2922
rect 27095 2922 33094 2950
rect 27095 -2922 33010 2922
rect 33074 -2922 33094 2922
rect 27095 -2950 33094 -2922
rect 33114 2922 39113 2950
rect 33114 -2922 39029 2922
rect 39093 -2922 39113 2922
rect 33114 -2950 39113 -2922
rect 39133 2922 45132 2950
rect 39133 -2922 45048 2922
rect 45112 -2922 45132 2922
rect 39133 -2950 45132 -2922
rect -45133 -3078 -39134 -3050
rect -45133 -8922 -39218 -3078
rect -39154 -8922 -39134 -3078
rect -45133 -8950 -39134 -8922
rect -39114 -3078 -33115 -3050
rect -39114 -8922 -33199 -3078
rect -33135 -8922 -33115 -3078
rect -39114 -8950 -33115 -8922
rect -33095 -3078 -27096 -3050
rect -33095 -8922 -27180 -3078
rect -27116 -8922 -27096 -3078
rect -33095 -8950 -27096 -8922
rect -27076 -3078 -21077 -3050
rect -27076 -8922 -21161 -3078
rect -21097 -8922 -21077 -3078
rect -27076 -8950 -21077 -8922
rect -21057 -3078 -15058 -3050
rect -21057 -8922 -15142 -3078
rect -15078 -8922 -15058 -3078
rect -21057 -8950 -15058 -8922
rect -15038 -3078 -9039 -3050
rect -15038 -8922 -9123 -3078
rect -9059 -8922 -9039 -3078
rect -15038 -8950 -9039 -8922
rect -9019 -3078 -3020 -3050
rect -9019 -8922 -3104 -3078
rect -3040 -8922 -3020 -3078
rect -9019 -8950 -3020 -8922
rect -3000 -3078 2999 -3050
rect -3000 -8922 2915 -3078
rect 2979 -8922 2999 -3078
rect -3000 -8950 2999 -8922
rect 3019 -3078 9018 -3050
rect 3019 -8922 8934 -3078
rect 8998 -8922 9018 -3078
rect 3019 -8950 9018 -8922
rect 9038 -3078 15037 -3050
rect 9038 -8922 14953 -3078
rect 15017 -8922 15037 -3078
rect 9038 -8950 15037 -8922
rect 15057 -3078 21056 -3050
rect 15057 -8922 20972 -3078
rect 21036 -8922 21056 -3078
rect 15057 -8950 21056 -8922
rect 21076 -3078 27075 -3050
rect 21076 -8922 26991 -3078
rect 27055 -8922 27075 -3078
rect 21076 -8950 27075 -8922
rect 27095 -3078 33094 -3050
rect 27095 -8922 33010 -3078
rect 33074 -8922 33094 -3078
rect 27095 -8950 33094 -8922
rect 33114 -3078 39113 -3050
rect 33114 -8922 39029 -3078
rect 39093 -8922 39113 -3078
rect 33114 -8950 39113 -8922
rect 39133 -3078 45132 -3050
rect 39133 -8922 45048 -3078
rect 45112 -8922 45132 -3078
rect 39133 -8950 45132 -8922
rect -45133 -9078 -39134 -9050
rect -45133 -14922 -39218 -9078
rect -39154 -14922 -39134 -9078
rect -45133 -14950 -39134 -14922
rect -39114 -9078 -33115 -9050
rect -39114 -14922 -33199 -9078
rect -33135 -14922 -33115 -9078
rect -39114 -14950 -33115 -14922
rect -33095 -9078 -27096 -9050
rect -33095 -14922 -27180 -9078
rect -27116 -14922 -27096 -9078
rect -33095 -14950 -27096 -14922
rect -27076 -9078 -21077 -9050
rect -27076 -14922 -21161 -9078
rect -21097 -14922 -21077 -9078
rect -27076 -14950 -21077 -14922
rect -21057 -9078 -15058 -9050
rect -21057 -14922 -15142 -9078
rect -15078 -14922 -15058 -9078
rect -21057 -14950 -15058 -14922
rect -15038 -9078 -9039 -9050
rect -15038 -14922 -9123 -9078
rect -9059 -14922 -9039 -9078
rect -15038 -14950 -9039 -14922
rect -9019 -9078 -3020 -9050
rect -9019 -14922 -3104 -9078
rect -3040 -14922 -3020 -9078
rect -9019 -14950 -3020 -14922
rect -3000 -9078 2999 -9050
rect -3000 -14922 2915 -9078
rect 2979 -14922 2999 -9078
rect -3000 -14950 2999 -14922
rect 3019 -9078 9018 -9050
rect 3019 -14922 8934 -9078
rect 8998 -14922 9018 -9078
rect 3019 -14950 9018 -14922
rect 9038 -9078 15037 -9050
rect 9038 -14922 14953 -9078
rect 15017 -14922 15037 -9078
rect 9038 -14950 15037 -14922
rect 15057 -9078 21056 -9050
rect 15057 -14922 20972 -9078
rect 21036 -14922 21056 -9078
rect 15057 -14950 21056 -14922
rect 21076 -9078 27075 -9050
rect 21076 -14922 26991 -9078
rect 27055 -14922 27075 -9078
rect 21076 -14950 27075 -14922
rect 27095 -9078 33094 -9050
rect 27095 -14922 33010 -9078
rect 33074 -14922 33094 -9078
rect 27095 -14950 33094 -14922
rect 33114 -9078 39113 -9050
rect 33114 -14922 39029 -9078
rect 39093 -14922 39113 -9078
rect 33114 -14950 39113 -14922
rect 39133 -9078 45132 -9050
rect 39133 -14922 45048 -9078
rect 45112 -14922 45132 -9078
rect 39133 -14950 45132 -14922
rect -45133 -15078 -39134 -15050
rect -45133 -20922 -39218 -15078
rect -39154 -20922 -39134 -15078
rect -45133 -20950 -39134 -20922
rect -39114 -15078 -33115 -15050
rect -39114 -20922 -33199 -15078
rect -33135 -20922 -33115 -15078
rect -39114 -20950 -33115 -20922
rect -33095 -15078 -27096 -15050
rect -33095 -20922 -27180 -15078
rect -27116 -20922 -27096 -15078
rect -33095 -20950 -27096 -20922
rect -27076 -15078 -21077 -15050
rect -27076 -20922 -21161 -15078
rect -21097 -20922 -21077 -15078
rect -27076 -20950 -21077 -20922
rect -21057 -15078 -15058 -15050
rect -21057 -20922 -15142 -15078
rect -15078 -20922 -15058 -15078
rect -21057 -20950 -15058 -20922
rect -15038 -15078 -9039 -15050
rect -15038 -20922 -9123 -15078
rect -9059 -20922 -9039 -15078
rect -15038 -20950 -9039 -20922
rect -9019 -15078 -3020 -15050
rect -9019 -20922 -3104 -15078
rect -3040 -20922 -3020 -15078
rect -9019 -20950 -3020 -20922
rect -3000 -15078 2999 -15050
rect -3000 -20922 2915 -15078
rect 2979 -20922 2999 -15078
rect -3000 -20950 2999 -20922
rect 3019 -15078 9018 -15050
rect 3019 -20922 8934 -15078
rect 8998 -20922 9018 -15078
rect 3019 -20950 9018 -20922
rect 9038 -15078 15037 -15050
rect 9038 -20922 14953 -15078
rect 15017 -20922 15037 -15078
rect 9038 -20950 15037 -20922
rect 15057 -15078 21056 -15050
rect 15057 -20922 20972 -15078
rect 21036 -20922 21056 -15078
rect 15057 -20950 21056 -20922
rect 21076 -15078 27075 -15050
rect 21076 -20922 26991 -15078
rect 27055 -20922 27075 -15078
rect 21076 -20950 27075 -20922
rect 27095 -15078 33094 -15050
rect 27095 -20922 33010 -15078
rect 33074 -20922 33094 -15078
rect 27095 -20950 33094 -20922
rect 33114 -15078 39113 -15050
rect 33114 -20922 39029 -15078
rect 39093 -20922 39113 -15078
rect 33114 -20950 39113 -20922
rect 39133 -15078 45132 -15050
rect 39133 -20922 45048 -15078
rect 45112 -20922 45132 -15078
rect 39133 -20950 45132 -20922
<< via3 >>
rect -39218 15078 -39154 20922
rect -33199 15078 -33135 20922
rect -27180 15078 -27116 20922
rect -21161 15078 -21097 20922
rect -15142 15078 -15078 20922
rect -9123 15078 -9059 20922
rect -3104 15078 -3040 20922
rect 2915 15078 2979 20922
rect 8934 15078 8998 20922
rect 14953 15078 15017 20922
rect 20972 15078 21036 20922
rect 26991 15078 27055 20922
rect 33010 15078 33074 20922
rect 39029 15078 39093 20922
rect 45048 15078 45112 20922
rect -39218 9078 -39154 14922
rect -33199 9078 -33135 14922
rect -27180 9078 -27116 14922
rect -21161 9078 -21097 14922
rect -15142 9078 -15078 14922
rect -9123 9078 -9059 14922
rect -3104 9078 -3040 14922
rect 2915 9078 2979 14922
rect 8934 9078 8998 14922
rect 14953 9078 15017 14922
rect 20972 9078 21036 14922
rect 26991 9078 27055 14922
rect 33010 9078 33074 14922
rect 39029 9078 39093 14922
rect 45048 9078 45112 14922
rect -39218 3078 -39154 8922
rect -33199 3078 -33135 8922
rect -27180 3078 -27116 8922
rect -21161 3078 -21097 8922
rect -15142 3078 -15078 8922
rect -9123 3078 -9059 8922
rect -3104 3078 -3040 8922
rect 2915 3078 2979 8922
rect 8934 3078 8998 8922
rect 14953 3078 15017 8922
rect 20972 3078 21036 8922
rect 26991 3078 27055 8922
rect 33010 3078 33074 8922
rect 39029 3078 39093 8922
rect 45048 3078 45112 8922
rect -39218 -2922 -39154 2922
rect -33199 -2922 -33135 2922
rect -27180 -2922 -27116 2922
rect -21161 -2922 -21097 2922
rect -15142 -2922 -15078 2922
rect -9123 -2922 -9059 2922
rect -3104 -2922 -3040 2922
rect 2915 -2922 2979 2922
rect 8934 -2922 8998 2922
rect 14953 -2922 15017 2922
rect 20972 -2922 21036 2922
rect 26991 -2922 27055 2922
rect 33010 -2922 33074 2922
rect 39029 -2922 39093 2922
rect 45048 -2922 45112 2922
rect -39218 -8922 -39154 -3078
rect -33199 -8922 -33135 -3078
rect -27180 -8922 -27116 -3078
rect -21161 -8922 -21097 -3078
rect -15142 -8922 -15078 -3078
rect -9123 -8922 -9059 -3078
rect -3104 -8922 -3040 -3078
rect 2915 -8922 2979 -3078
rect 8934 -8922 8998 -3078
rect 14953 -8922 15017 -3078
rect 20972 -8922 21036 -3078
rect 26991 -8922 27055 -3078
rect 33010 -8922 33074 -3078
rect 39029 -8922 39093 -3078
rect 45048 -8922 45112 -3078
rect -39218 -14922 -39154 -9078
rect -33199 -14922 -33135 -9078
rect -27180 -14922 -27116 -9078
rect -21161 -14922 -21097 -9078
rect -15142 -14922 -15078 -9078
rect -9123 -14922 -9059 -9078
rect -3104 -14922 -3040 -9078
rect 2915 -14922 2979 -9078
rect 8934 -14922 8998 -9078
rect 14953 -14922 15017 -9078
rect 20972 -14922 21036 -9078
rect 26991 -14922 27055 -9078
rect 33010 -14922 33074 -9078
rect 39029 -14922 39093 -9078
rect 45048 -14922 45112 -9078
rect -39218 -20922 -39154 -15078
rect -33199 -20922 -33135 -15078
rect -27180 -20922 -27116 -15078
rect -21161 -20922 -21097 -15078
rect -15142 -20922 -15078 -15078
rect -9123 -20922 -9059 -15078
rect -3104 -20922 -3040 -15078
rect 2915 -20922 2979 -15078
rect 8934 -20922 8998 -15078
rect 14953 -20922 15017 -15078
rect 20972 -20922 21036 -15078
rect 26991 -20922 27055 -15078
rect 33010 -20922 33074 -15078
rect 39029 -20922 39093 -15078
rect 45048 -20922 45112 -15078
<< mimcap >>
rect -45033 20810 -39333 20850
rect -45033 15190 -44993 20810
rect -39373 15190 -39333 20810
rect -45033 15150 -39333 15190
rect -39014 20810 -33314 20850
rect -39014 15190 -38974 20810
rect -33354 15190 -33314 20810
rect -39014 15150 -33314 15190
rect -32995 20810 -27295 20850
rect -32995 15190 -32955 20810
rect -27335 15190 -27295 20810
rect -32995 15150 -27295 15190
rect -26976 20810 -21276 20850
rect -26976 15190 -26936 20810
rect -21316 15190 -21276 20810
rect -26976 15150 -21276 15190
rect -20957 20810 -15257 20850
rect -20957 15190 -20917 20810
rect -15297 15190 -15257 20810
rect -20957 15150 -15257 15190
rect -14938 20810 -9238 20850
rect -14938 15190 -14898 20810
rect -9278 15190 -9238 20810
rect -14938 15150 -9238 15190
rect -8919 20810 -3219 20850
rect -8919 15190 -8879 20810
rect -3259 15190 -3219 20810
rect -8919 15150 -3219 15190
rect -2900 20810 2800 20850
rect -2900 15190 -2860 20810
rect 2760 15190 2800 20810
rect -2900 15150 2800 15190
rect 3119 20810 8819 20850
rect 3119 15190 3159 20810
rect 8779 15190 8819 20810
rect 3119 15150 8819 15190
rect 9138 20810 14838 20850
rect 9138 15190 9178 20810
rect 14798 15190 14838 20810
rect 9138 15150 14838 15190
rect 15157 20810 20857 20850
rect 15157 15190 15197 20810
rect 20817 15190 20857 20810
rect 15157 15150 20857 15190
rect 21176 20810 26876 20850
rect 21176 15190 21216 20810
rect 26836 15190 26876 20810
rect 21176 15150 26876 15190
rect 27195 20810 32895 20850
rect 27195 15190 27235 20810
rect 32855 15190 32895 20810
rect 27195 15150 32895 15190
rect 33214 20810 38914 20850
rect 33214 15190 33254 20810
rect 38874 15190 38914 20810
rect 33214 15150 38914 15190
rect 39233 20810 44933 20850
rect 39233 15190 39273 20810
rect 44893 15190 44933 20810
rect 39233 15150 44933 15190
rect -45033 14810 -39333 14850
rect -45033 9190 -44993 14810
rect -39373 9190 -39333 14810
rect -45033 9150 -39333 9190
rect -39014 14810 -33314 14850
rect -39014 9190 -38974 14810
rect -33354 9190 -33314 14810
rect -39014 9150 -33314 9190
rect -32995 14810 -27295 14850
rect -32995 9190 -32955 14810
rect -27335 9190 -27295 14810
rect -32995 9150 -27295 9190
rect -26976 14810 -21276 14850
rect -26976 9190 -26936 14810
rect -21316 9190 -21276 14810
rect -26976 9150 -21276 9190
rect -20957 14810 -15257 14850
rect -20957 9190 -20917 14810
rect -15297 9190 -15257 14810
rect -20957 9150 -15257 9190
rect -14938 14810 -9238 14850
rect -14938 9190 -14898 14810
rect -9278 9190 -9238 14810
rect -14938 9150 -9238 9190
rect -8919 14810 -3219 14850
rect -8919 9190 -8879 14810
rect -3259 9190 -3219 14810
rect -8919 9150 -3219 9190
rect -2900 14810 2800 14850
rect -2900 9190 -2860 14810
rect 2760 9190 2800 14810
rect -2900 9150 2800 9190
rect 3119 14810 8819 14850
rect 3119 9190 3159 14810
rect 8779 9190 8819 14810
rect 3119 9150 8819 9190
rect 9138 14810 14838 14850
rect 9138 9190 9178 14810
rect 14798 9190 14838 14810
rect 9138 9150 14838 9190
rect 15157 14810 20857 14850
rect 15157 9190 15197 14810
rect 20817 9190 20857 14810
rect 15157 9150 20857 9190
rect 21176 14810 26876 14850
rect 21176 9190 21216 14810
rect 26836 9190 26876 14810
rect 21176 9150 26876 9190
rect 27195 14810 32895 14850
rect 27195 9190 27235 14810
rect 32855 9190 32895 14810
rect 27195 9150 32895 9190
rect 33214 14810 38914 14850
rect 33214 9190 33254 14810
rect 38874 9190 38914 14810
rect 33214 9150 38914 9190
rect 39233 14810 44933 14850
rect 39233 9190 39273 14810
rect 44893 9190 44933 14810
rect 39233 9150 44933 9190
rect -45033 8810 -39333 8850
rect -45033 3190 -44993 8810
rect -39373 3190 -39333 8810
rect -45033 3150 -39333 3190
rect -39014 8810 -33314 8850
rect -39014 3190 -38974 8810
rect -33354 3190 -33314 8810
rect -39014 3150 -33314 3190
rect -32995 8810 -27295 8850
rect -32995 3190 -32955 8810
rect -27335 3190 -27295 8810
rect -32995 3150 -27295 3190
rect -26976 8810 -21276 8850
rect -26976 3190 -26936 8810
rect -21316 3190 -21276 8810
rect -26976 3150 -21276 3190
rect -20957 8810 -15257 8850
rect -20957 3190 -20917 8810
rect -15297 3190 -15257 8810
rect -20957 3150 -15257 3190
rect -14938 8810 -9238 8850
rect -14938 3190 -14898 8810
rect -9278 3190 -9238 8810
rect -14938 3150 -9238 3190
rect -8919 8810 -3219 8850
rect -8919 3190 -8879 8810
rect -3259 3190 -3219 8810
rect -8919 3150 -3219 3190
rect -2900 8810 2800 8850
rect -2900 3190 -2860 8810
rect 2760 3190 2800 8810
rect -2900 3150 2800 3190
rect 3119 8810 8819 8850
rect 3119 3190 3159 8810
rect 8779 3190 8819 8810
rect 3119 3150 8819 3190
rect 9138 8810 14838 8850
rect 9138 3190 9178 8810
rect 14798 3190 14838 8810
rect 9138 3150 14838 3190
rect 15157 8810 20857 8850
rect 15157 3190 15197 8810
rect 20817 3190 20857 8810
rect 15157 3150 20857 3190
rect 21176 8810 26876 8850
rect 21176 3190 21216 8810
rect 26836 3190 26876 8810
rect 21176 3150 26876 3190
rect 27195 8810 32895 8850
rect 27195 3190 27235 8810
rect 32855 3190 32895 8810
rect 27195 3150 32895 3190
rect 33214 8810 38914 8850
rect 33214 3190 33254 8810
rect 38874 3190 38914 8810
rect 33214 3150 38914 3190
rect 39233 8810 44933 8850
rect 39233 3190 39273 8810
rect 44893 3190 44933 8810
rect 39233 3150 44933 3190
rect -45033 2810 -39333 2850
rect -45033 -2810 -44993 2810
rect -39373 -2810 -39333 2810
rect -45033 -2850 -39333 -2810
rect -39014 2810 -33314 2850
rect -39014 -2810 -38974 2810
rect -33354 -2810 -33314 2810
rect -39014 -2850 -33314 -2810
rect -32995 2810 -27295 2850
rect -32995 -2810 -32955 2810
rect -27335 -2810 -27295 2810
rect -32995 -2850 -27295 -2810
rect -26976 2810 -21276 2850
rect -26976 -2810 -26936 2810
rect -21316 -2810 -21276 2810
rect -26976 -2850 -21276 -2810
rect -20957 2810 -15257 2850
rect -20957 -2810 -20917 2810
rect -15297 -2810 -15257 2810
rect -20957 -2850 -15257 -2810
rect -14938 2810 -9238 2850
rect -14938 -2810 -14898 2810
rect -9278 -2810 -9238 2810
rect -14938 -2850 -9238 -2810
rect -8919 2810 -3219 2850
rect -8919 -2810 -8879 2810
rect -3259 -2810 -3219 2810
rect -8919 -2850 -3219 -2810
rect -2900 2810 2800 2850
rect -2900 -2810 -2860 2810
rect 2760 -2810 2800 2810
rect -2900 -2850 2800 -2810
rect 3119 2810 8819 2850
rect 3119 -2810 3159 2810
rect 8779 -2810 8819 2810
rect 3119 -2850 8819 -2810
rect 9138 2810 14838 2850
rect 9138 -2810 9178 2810
rect 14798 -2810 14838 2810
rect 9138 -2850 14838 -2810
rect 15157 2810 20857 2850
rect 15157 -2810 15197 2810
rect 20817 -2810 20857 2810
rect 15157 -2850 20857 -2810
rect 21176 2810 26876 2850
rect 21176 -2810 21216 2810
rect 26836 -2810 26876 2810
rect 21176 -2850 26876 -2810
rect 27195 2810 32895 2850
rect 27195 -2810 27235 2810
rect 32855 -2810 32895 2810
rect 27195 -2850 32895 -2810
rect 33214 2810 38914 2850
rect 33214 -2810 33254 2810
rect 38874 -2810 38914 2810
rect 33214 -2850 38914 -2810
rect 39233 2810 44933 2850
rect 39233 -2810 39273 2810
rect 44893 -2810 44933 2810
rect 39233 -2850 44933 -2810
rect -45033 -3190 -39333 -3150
rect -45033 -8810 -44993 -3190
rect -39373 -8810 -39333 -3190
rect -45033 -8850 -39333 -8810
rect -39014 -3190 -33314 -3150
rect -39014 -8810 -38974 -3190
rect -33354 -8810 -33314 -3190
rect -39014 -8850 -33314 -8810
rect -32995 -3190 -27295 -3150
rect -32995 -8810 -32955 -3190
rect -27335 -8810 -27295 -3190
rect -32995 -8850 -27295 -8810
rect -26976 -3190 -21276 -3150
rect -26976 -8810 -26936 -3190
rect -21316 -8810 -21276 -3190
rect -26976 -8850 -21276 -8810
rect -20957 -3190 -15257 -3150
rect -20957 -8810 -20917 -3190
rect -15297 -8810 -15257 -3190
rect -20957 -8850 -15257 -8810
rect -14938 -3190 -9238 -3150
rect -14938 -8810 -14898 -3190
rect -9278 -8810 -9238 -3190
rect -14938 -8850 -9238 -8810
rect -8919 -3190 -3219 -3150
rect -8919 -8810 -8879 -3190
rect -3259 -8810 -3219 -3190
rect -8919 -8850 -3219 -8810
rect -2900 -3190 2800 -3150
rect -2900 -8810 -2860 -3190
rect 2760 -8810 2800 -3190
rect -2900 -8850 2800 -8810
rect 3119 -3190 8819 -3150
rect 3119 -8810 3159 -3190
rect 8779 -8810 8819 -3190
rect 3119 -8850 8819 -8810
rect 9138 -3190 14838 -3150
rect 9138 -8810 9178 -3190
rect 14798 -8810 14838 -3190
rect 9138 -8850 14838 -8810
rect 15157 -3190 20857 -3150
rect 15157 -8810 15197 -3190
rect 20817 -8810 20857 -3190
rect 15157 -8850 20857 -8810
rect 21176 -3190 26876 -3150
rect 21176 -8810 21216 -3190
rect 26836 -8810 26876 -3190
rect 21176 -8850 26876 -8810
rect 27195 -3190 32895 -3150
rect 27195 -8810 27235 -3190
rect 32855 -8810 32895 -3190
rect 27195 -8850 32895 -8810
rect 33214 -3190 38914 -3150
rect 33214 -8810 33254 -3190
rect 38874 -8810 38914 -3190
rect 33214 -8850 38914 -8810
rect 39233 -3190 44933 -3150
rect 39233 -8810 39273 -3190
rect 44893 -8810 44933 -3190
rect 39233 -8850 44933 -8810
rect -45033 -9190 -39333 -9150
rect -45033 -14810 -44993 -9190
rect -39373 -14810 -39333 -9190
rect -45033 -14850 -39333 -14810
rect -39014 -9190 -33314 -9150
rect -39014 -14810 -38974 -9190
rect -33354 -14810 -33314 -9190
rect -39014 -14850 -33314 -14810
rect -32995 -9190 -27295 -9150
rect -32995 -14810 -32955 -9190
rect -27335 -14810 -27295 -9190
rect -32995 -14850 -27295 -14810
rect -26976 -9190 -21276 -9150
rect -26976 -14810 -26936 -9190
rect -21316 -14810 -21276 -9190
rect -26976 -14850 -21276 -14810
rect -20957 -9190 -15257 -9150
rect -20957 -14810 -20917 -9190
rect -15297 -14810 -15257 -9190
rect -20957 -14850 -15257 -14810
rect -14938 -9190 -9238 -9150
rect -14938 -14810 -14898 -9190
rect -9278 -14810 -9238 -9190
rect -14938 -14850 -9238 -14810
rect -8919 -9190 -3219 -9150
rect -8919 -14810 -8879 -9190
rect -3259 -14810 -3219 -9190
rect -8919 -14850 -3219 -14810
rect -2900 -9190 2800 -9150
rect -2900 -14810 -2860 -9190
rect 2760 -14810 2800 -9190
rect -2900 -14850 2800 -14810
rect 3119 -9190 8819 -9150
rect 3119 -14810 3159 -9190
rect 8779 -14810 8819 -9190
rect 3119 -14850 8819 -14810
rect 9138 -9190 14838 -9150
rect 9138 -14810 9178 -9190
rect 14798 -14810 14838 -9190
rect 9138 -14850 14838 -14810
rect 15157 -9190 20857 -9150
rect 15157 -14810 15197 -9190
rect 20817 -14810 20857 -9190
rect 15157 -14850 20857 -14810
rect 21176 -9190 26876 -9150
rect 21176 -14810 21216 -9190
rect 26836 -14810 26876 -9190
rect 21176 -14850 26876 -14810
rect 27195 -9190 32895 -9150
rect 27195 -14810 27235 -9190
rect 32855 -14810 32895 -9190
rect 27195 -14850 32895 -14810
rect 33214 -9190 38914 -9150
rect 33214 -14810 33254 -9190
rect 38874 -14810 38914 -9190
rect 33214 -14850 38914 -14810
rect 39233 -9190 44933 -9150
rect 39233 -14810 39273 -9190
rect 44893 -14810 44933 -9190
rect 39233 -14850 44933 -14810
rect -45033 -15190 -39333 -15150
rect -45033 -20810 -44993 -15190
rect -39373 -20810 -39333 -15190
rect -45033 -20850 -39333 -20810
rect -39014 -15190 -33314 -15150
rect -39014 -20810 -38974 -15190
rect -33354 -20810 -33314 -15190
rect -39014 -20850 -33314 -20810
rect -32995 -15190 -27295 -15150
rect -32995 -20810 -32955 -15190
rect -27335 -20810 -27295 -15190
rect -32995 -20850 -27295 -20810
rect -26976 -15190 -21276 -15150
rect -26976 -20810 -26936 -15190
rect -21316 -20810 -21276 -15190
rect -26976 -20850 -21276 -20810
rect -20957 -15190 -15257 -15150
rect -20957 -20810 -20917 -15190
rect -15297 -20810 -15257 -15190
rect -20957 -20850 -15257 -20810
rect -14938 -15190 -9238 -15150
rect -14938 -20810 -14898 -15190
rect -9278 -20810 -9238 -15190
rect -14938 -20850 -9238 -20810
rect -8919 -15190 -3219 -15150
rect -8919 -20810 -8879 -15190
rect -3259 -20810 -3219 -15190
rect -8919 -20850 -3219 -20810
rect -2900 -15190 2800 -15150
rect -2900 -20810 -2860 -15190
rect 2760 -20810 2800 -15190
rect -2900 -20850 2800 -20810
rect 3119 -15190 8819 -15150
rect 3119 -20810 3159 -15190
rect 8779 -20810 8819 -15190
rect 3119 -20850 8819 -20810
rect 9138 -15190 14838 -15150
rect 9138 -20810 9178 -15190
rect 14798 -20810 14838 -15190
rect 9138 -20850 14838 -20810
rect 15157 -15190 20857 -15150
rect 15157 -20810 15197 -15190
rect 20817 -20810 20857 -15190
rect 15157 -20850 20857 -20810
rect 21176 -15190 26876 -15150
rect 21176 -20810 21216 -15190
rect 26836 -20810 26876 -15190
rect 21176 -20850 26876 -20810
rect 27195 -15190 32895 -15150
rect 27195 -20810 27235 -15190
rect 32855 -20810 32895 -15190
rect 27195 -20850 32895 -20810
rect 33214 -15190 38914 -15150
rect 33214 -20810 33254 -15190
rect 38874 -20810 38914 -15190
rect 33214 -20850 38914 -20810
rect 39233 -15190 44933 -15150
rect 39233 -20810 39273 -15190
rect 44893 -20810 44933 -15190
rect 39233 -20850 44933 -20810
<< mimcapcontact >>
rect -44993 15190 -39373 20810
rect -38974 15190 -33354 20810
rect -32955 15190 -27335 20810
rect -26936 15190 -21316 20810
rect -20917 15190 -15297 20810
rect -14898 15190 -9278 20810
rect -8879 15190 -3259 20810
rect -2860 15190 2760 20810
rect 3159 15190 8779 20810
rect 9178 15190 14798 20810
rect 15197 15190 20817 20810
rect 21216 15190 26836 20810
rect 27235 15190 32855 20810
rect 33254 15190 38874 20810
rect 39273 15190 44893 20810
rect -44993 9190 -39373 14810
rect -38974 9190 -33354 14810
rect -32955 9190 -27335 14810
rect -26936 9190 -21316 14810
rect -20917 9190 -15297 14810
rect -14898 9190 -9278 14810
rect -8879 9190 -3259 14810
rect -2860 9190 2760 14810
rect 3159 9190 8779 14810
rect 9178 9190 14798 14810
rect 15197 9190 20817 14810
rect 21216 9190 26836 14810
rect 27235 9190 32855 14810
rect 33254 9190 38874 14810
rect 39273 9190 44893 14810
rect -44993 3190 -39373 8810
rect -38974 3190 -33354 8810
rect -32955 3190 -27335 8810
rect -26936 3190 -21316 8810
rect -20917 3190 -15297 8810
rect -14898 3190 -9278 8810
rect -8879 3190 -3259 8810
rect -2860 3190 2760 8810
rect 3159 3190 8779 8810
rect 9178 3190 14798 8810
rect 15197 3190 20817 8810
rect 21216 3190 26836 8810
rect 27235 3190 32855 8810
rect 33254 3190 38874 8810
rect 39273 3190 44893 8810
rect -44993 -2810 -39373 2810
rect -38974 -2810 -33354 2810
rect -32955 -2810 -27335 2810
rect -26936 -2810 -21316 2810
rect -20917 -2810 -15297 2810
rect -14898 -2810 -9278 2810
rect -8879 -2810 -3259 2810
rect -2860 -2810 2760 2810
rect 3159 -2810 8779 2810
rect 9178 -2810 14798 2810
rect 15197 -2810 20817 2810
rect 21216 -2810 26836 2810
rect 27235 -2810 32855 2810
rect 33254 -2810 38874 2810
rect 39273 -2810 44893 2810
rect -44993 -8810 -39373 -3190
rect -38974 -8810 -33354 -3190
rect -32955 -8810 -27335 -3190
rect -26936 -8810 -21316 -3190
rect -20917 -8810 -15297 -3190
rect -14898 -8810 -9278 -3190
rect -8879 -8810 -3259 -3190
rect -2860 -8810 2760 -3190
rect 3159 -8810 8779 -3190
rect 9178 -8810 14798 -3190
rect 15197 -8810 20817 -3190
rect 21216 -8810 26836 -3190
rect 27235 -8810 32855 -3190
rect 33254 -8810 38874 -3190
rect 39273 -8810 44893 -3190
rect -44993 -14810 -39373 -9190
rect -38974 -14810 -33354 -9190
rect -32955 -14810 -27335 -9190
rect -26936 -14810 -21316 -9190
rect -20917 -14810 -15297 -9190
rect -14898 -14810 -9278 -9190
rect -8879 -14810 -3259 -9190
rect -2860 -14810 2760 -9190
rect 3159 -14810 8779 -9190
rect 9178 -14810 14798 -9190
rect 15197 -14810 20817 -9190
rect 21216 -14810 26836 -9190
rect 27235 -14810 32855 -9190
rect 33254 -14810 38874 -9190
rect 39273 -14810 44893 -9190
rect -44993 -20810 -39373 -15190
rect -38974 -20810 -33354 -15190
rect -32955 -20810 -27335 -15190
rect -26936 -20810 -21316 -15190
rect -20917 -20810 -15297 -15190
rect -14898 -20810 -9278 -15190
rect -8879 -20810 -3259 -15190
rect -2860 -20810 2760 -15190
rect 3159 -20810 8779 -15190
rect 9178 -20810 14798 -15190
rect 15197 -20810 20817 -15190
rect 21216 -20810 26836 -15190
rect 27235 -20810 32855 -15190
rect 33254 -20810 38874 -15190
rect 39273 -20810 44893 -15190
<< metal4 >>
rect -39265 20938 -39161 21000
rect -33246 20938 -33142 21000
rect -27227 20938 -27123 21000
rect -21208 20938 -21104 21000
rect -15189 20938 -15085 21000
rect -9170 20938 -9066 21000
rect -3151 20938 -3047 21000
rect 2868 20938 2972 21000
rect 8887 20938 8991 21000
rect 14906 20938 15010 21000
rect 20925 20938 21029 21000
rect 26944 20938 27048 21000
rect 32963 20938 33067 21000
rect 38982 20938 39086 21000
rect 45001 20938 45105 21000
rect -39265 20922 -39138 20938
rect -44994 20810 -39372 20811
rect -44994 15190 -44993 20810
rect -39373 15190 -39372 20810
rect -44994 15189 -39372 15190
rect -39265 15078 -39218 20922
rect -39154 15078 -39138 20922
rect -33246 20922 -33119 20938
rect -38975 20810 -33353 20811
rect -38975 15190 -38974 20810
rect -33354 15190 -33353 20810
rect -38975 15189 -33353 15190
rect -39265 15062 -39138 15078
rect -33246 15078 -33199 20922
rect -33135 15078 -33119 20922
rect -27227 20922 -27100 20938
rect -32956 20810 -27334 20811
rect -32956 15190 -32955 20810
rect -27335 15190 -27334 20810
rect -32956 15189 -27334 15190
rect -33246 15062 -33119 15078
rect -27227 15078 -27180 20922
rect -27116 15078 -27100 20922
rect -21208 20922 -21081 20938
rect -26937 20810 -21315 20811
rect -26937 15190 -26936 20810
rect -21316 15190 -21315 20810
rect -26937 15189 -21315 15190
rect -27227 15062 -27100 15078
rect -21208 15078 -21161 20922
rect -21097 15078 -21081 20922
rect -15189 20922 -15062 20938
rect -20918 20810 -15296 20811
rect -20918 15190 -20917 20810
rect -15297 15190 -15296 20810
rect -20918 15189 -15296 15190
rect -21208 15062 -21081 15078
rect -15189 15078 -15142 20922
rect -15078 15078 -15062 20922
rect -9170 20922 -9043 20938
rect -14899 20810 -9277 20811
rect -14899 15190 -14898 20810
rect -9278 15190 -9277 20810
rect -14899 15189 -9277 15190
rect -15189 15062 -15062 15078
rect -9170 15078 -9123 20922
rect -9059 15078 -9043 20922
rect -3151 20922 -3024 20938
rect -8880 20810 -3258 20811
rect -8880 15190 -8879 20810
rect -3259 15190 -3258 20810
rect -8880 15189 -3258 15190
rect -9170 15062 -9043 15078
rect -3151 15078 -3104 20922
rect -3040 15078 -3024 20922
rect 2868 20922 2995 20938
rect -2861 20810 2761 20811
rect -2861 15190 -2860 20810
rect 2760 15190 2761 20810
rect -2861 15189 2761 15190
rect -3151 15062 -3024 15078
rect 2868 15078 2915 20922
rect 2979 15078 2995 20922
rect 8887 20922 9014 20938
rect 3158 20810 8780 20811
rect 3158 15190 3159 20810
rect 8779 15190 8780 20810
rect 3158 15189 8780 15190
rect 2868 15062 2995 15078
rect 8887 15078 8934 20922
rect 8998 15078 9014 20922
rect 14906 20922 15033 20938
rect 9177 20810 14799 20811
rect 9177 15190 9178 20810
rect 14798 15190 14799 20810
rect 9177 15189 14799 15190
rect 8887 15062 9014 15078
rect 14906 15078 14953 20922
rect 15017 15078 15033 20922
rect 20925 20922 21052 20938
rect 15196 20810 20818 20811
rect 15196 15190 15197 20810
rect 20817 15190 20818 20810
rect 15196 15189 20818 15190
rect 14906 15062 15033 15078
rect 20925 15078 20972 20922
rect 21036 15078 21052 20922
rect 26944 20922 27071 20938
rect 21215 20810 26837 20811
rect 21215 15190 21216 20810
rect 26836 15190 26837 20810
rect 21215 15189 26837 15190
rect 20925 15062 21052 15078
rect 26944 15078 26991 20922
rect 27055 15078 27071 20922
rect 32963 20922 33090 20938
rect 27234 20810 32856 20811
rect 27234 15190 27235 20810
rect 32855 15190 32856 20810
rect 27234 15189 32856 15190
rect 26944 15062 27071 15078
rect 32963 15078 33010 20922
rect 33074 15078 33090 20922
rect 38982 20922 39109 20938
rect 33253 20810 38875 20811
rect 33253 15190 33254 20810
rect 38874 15190 38875 20810
rect 33253 15189 38875 15190
rect 32963 15062 33090 15078
rect 38982 15078 39029 20922
rect 39093 15078 39109 20922
rect 45001 20922 45128 20938
rect 39272 20810 44894 20811
rect 39272 15190 39273 20810
rect 44893 15190 44894 20810
rect 39272 15189 44894 15190
rect 38982 15062 39109 15078
rect 45001 15078 45048 20922
rect 45112 15078 45128 20922
rect 45001 15062 45128 15078
rect -39265 14938 -39161 15062
rect -33246 14938 -33142 15062
rect -27227 14938 -27123 15062
rect -21208 14938 -21104 15062
rect -15189 14938 -15085 15062
rect -9170 14938 -9066 15062
rect -3151 14938 -3047 15062
rect 2868 14938 2972 15062
rect 8887 14938 8991 15062
rect 14906 14938 15010 15062
rect 20925 14938 21029 15062
rect 26944 14938 27048 15062
rect 32963 14938 33067 15062
rect 38982 14938 39086 15062
rect 45001 14938 45105 15062
rect -39265 14922 -39138 14938
rect -44994 14810 -39372 14811
rect -44994 9190 -44993 14810
rect -39373 9190 -39372 14810
rect -44994 9189 -39372 9190
rect -39265 9078 -39218 14922
rect -39154 9078 -39138 14922
rect -33246 14922 -33119 14938
rect -38975 14810 -33353 14811
rect -38975 9190 -38974 14810
rect -33354 9190 -33353 14810
rect -38975 9189 -33353 9190
rect -39265 9062 -39138 9078
rect -33246 9078 -33199 14922
rect -33135 9078 -33119 14922
rect -27227 14922 -27100 14938
rect -32956 14810 -27334 14811
rect -32956 9190 -32955 14810
rect -27335 9190 -27334 14810
rect -32956 9189 -27334 9190
rect -33246 9062 -33119 9078
rect -27227 9078 -27180 14922
rect -27116 9078 -27100 14922
rect -21208 14922 -21081 14938
rect -26937 14810 -21315 14811
rect -26937 9190 -26936 14810
rect -21316 9190 -21315 14810
rect -26937 9189 -21315 9190
rect -27227 9062 -27100 9078
rect -21208 9078 -21161 14922
rect -21097 9078 -21081 14922
rect -15189 14922 -15062 14938
rect -20918 14810 -15296 14811
rect -20918 9190 -20917 14810
rect -15297 9190 -15296 14810
rect -20918 9189 -15296 9190
rect -21208 9062 -21081 9078
rect -15189 9078 -15142 14922
rect -15078 9078 -15062 14922
rect -9170 14922 -9043 14938
rect -14899 14810 -9277 14811
rect -14899 9190 -14898 14810
rect -9278 9190 -9277 14810
rect -14899 9189 -9277 9190
rect -15189 9062 -15062 9078
rect -9170 9078 -9123 14922
rect -9059 9078 -9043 14922
rect -3151 14922 -3024 14938
rect -8880 14810 -3258 14811
rect -8880 9190 -8879 14810
rect -3259 9190 -3258 14810
rect -8880 9189 -3258 9190
rect -9170 9062 -9043 9078
rect -3151 9078 -3104 14922
rect -3040 9078 -3024 14922
rect 2868 14922 2995 14938
rect -2861 14810 2761 14811
rect -2861 9190 -2860 14810
rect 2760 9190 2761 14810
rect -2861 9189 2761 9190
rect -3151 9062 -3024 9078
rect 2868 9078 2915 14922
rect 2979 9078 2995 14922
rect 8887 14922 9014 14938
rect 3158 14810 8780 14811
rect 3158 9190 3159 14810
rect 8779 9190 8780 14810
rect 3158 9189 8780 9190
rect 2868 9062 2995 9078
rect 8887 9078 8934 14922
rect 8998 9078 9014 14922
rect 14906 14922 15033 14938
rect 9177 14810 14799 14811
rect 9177 9190 9178 14810
rect 14798 9190 14799 14810
rect 9177 9189 14799 9190
rect 8887 9062 9014 9078
rect 14906 9078 14953 14922
rect 15017 9078 15033 14922
rect 20925 14922 21052 14938
rect 15196 14810 20818 14811
rect 15196 9190 15197 14810
rect 20817 9190 20818 14810
rect 15196 9189 20818 9190
rect 14906 9062 15033 9078
rect 20925 9078 20972 14922
rect 21036 9078 21052 14922
rect 26944 14922 27071 14938
rect 21215 14810 26837 14811
rect 21215 9190 21216 14810
rect 26836 9190 26837 14810
rect 21215 9189 26837 9190
rect 20925 9062 21052 9078
rect 26944 9078 26991 14922
rect 27055 9078 27071 14922
rect 32963 14922 33090 14938
rect 27234 14810 32856 14811
rect 27234 9190 27235 14810
rect 32855 9190 32856 14810
rect 27234 9189 32856 9190
rect 26944 9062 27071 9078
rect 32963 9078 33010 14922
rect 33074 9078 33090 14922
rect 38982 14922 39109 14938
rect 33253 14810 38875 14811
rect 33253 9190 33254 14810
rect 38874 9190 38875 14810
rect 33253 9189 38875 9190
rect 32963 9062 33090 9078
rect 38982 9078 39029 14922
rect 39093 9078 39109 14922
rect 45001 14922 45128 14938
rect 39272 14810 44894 14811
rect 39272 9190 39273 14810
rect 44893 9190 44894 14810
rect 39272 9189 44894 9190
rect 38982 9062 39109 9078
rect 45001 9078 45048 14922
rect 45112 9078 45128 14922
rect 45001 9062 45128 9078
rect -39265 8938 -39161 9062
rect -33246 8938 -33142 9062
rect -27227 8938 -27123 9062
rect -21208 8938 -21104 9062
rect -15189 8938 -15085 9062
rect -9170 8938 -9066 9062
rect -3151 8938 -3047 9062
rect 2868 8938 2972 9062
rect 8887 8938 8991 9062
rect 14906 8938 15010 9062
rect 20925 8938 21029 9062
rect 26944 8938 27048 9062
rect 32963 8938 33067 9062
rect 38982 8938 39086 9062
rect 45001 8938 45105 9062
rect -39265 8922 -39138 8938
rect -44994 8810 -39372 8811
rect -44994 3190 -44993 8810
rect -39373 3190 -39372 8810
rect -44994 3189 -39372 3190
rect -39265 3078 -39218 8922
rect -39154 3078 -39138 8922
rect -33246 8922 -33119 8938
rect -38975 8810 -33353 8811
rect -38975 3190 -38974 8810
rect -33354 3190 -33353 8810
rect -38975 3189 -33353 3190
rect -39265 3062 -39138 3078
rect -33246 3078 -33199 8922
rect -33135 3078 -33119 8922
rect -27227 8922 -27100 8938
rect -32956 8810 -27334 8811
rect -32956 3190 -32955 8810
rect -27335 3190 -27334 8810
rect -32956 3189 -27334 3190
rect -33246 3062 -33119 3078
rect -27227 3078 -27180 8922
rect -27116 3078 -27100 8922
rect -21208 8922 -21081 8938
rect -26937 8810 -21315 8811
rect -26937 3190 -26936 8810
rect -21316 3190 -21315 8810
rect -26937 3189 -21315 3190
rect -27227 3062 -27100 3078
rect -21208 3078 -21161 8922
rect -21097 3078 -21081 8922
rect -15189 8922 -15062 8938
rect -20918 8810 -15296 8811
rect -20918 3190 -20917 8810
rect -15297 3190 -15296 8810
rect -20918 3189 -15296 3190
rect -21208 3062 -21081 3078
rect -15189 3078 -15142 8922
rect -15078 3078 -15062 8922
rect -9170 8922 -9043 8938
rect -14899 8810 -9277 8811
rect -14899 3190 -14898 8810
rect -9278 3190 -9277 8810
rect -14899 3189 -9277 3190
rect -15189 3062 -15062 3078
rect -9170 3078 -9123 8922
rect -9059 3078 -9043 8922
rect -3151 8922 -3024 8938
rect -8880 8810 -3258 8811
rect -8880 3190 -8879 8810
rect -3259 3190 -3258 8810
rect -8880 3189 -3258 3190
rect -9170 3062 -9043 3078
rect -3151 3078 -3104 8922
rect -3040 3078 -3024 8922
rect 2868 8922 2995 8938
rect -2861 8810 2761 8811
rect -2861 3190 -2860 8810
rect 2760 3190 2761 8810
rect -2861 3189 2761 3190
rect -3151 3062 -3024 3078
rect 2868 3078 2915 8922
rect 2979 3078 2995 8922
rect 8887 8922 9014 8938
rect 3158 8810 8780 8811
rect 3158 3190 3159 8810
rect 8779 3190 8780 8810
rect 3158 3189 8780 3190
rect 2868 3062 2995 3078
rect 8887 3078 8934 8922
rect 8998 3078 9014 8922
rect 14906 8922 15033 8938
rect 9177 8810 14799 8811
rect 9177 3190 9178 8810
rect 14798 3190 14799 8810
rect 9177 3189 14799 3190
rect 8887 3062 9014 3078
rect 14906 3078 14953 8922
rect 15017 3078 15033 8922
rect 20925 8922 21052 8938
rect 15196 8810 20818 8811
rect 15196 3190 15197 8810
rect 20817 3190 20818 8810
rect 15196 3189 20818 3190
rect 14906 3062 15033 3078
rect 20925 3078 20972 8922
rect 21036 3078 21052 8922
rect 26944 8922 27071 8938
rect 21215 8810 26837 8811
rect 21215 3190 21216 8810
rect 26836 3190 26837 8810
rect 21215 3189 26837 3190
rect 20925 3062 21052 3078
rect 26944 3078 26991 8922
rect 27055 3078 27071 8922
rect 32963 8922 33090 8938
rect 27234 8810 32856 8811
rect 27234 3190 27235 8810
rect 32855 3190 32856 8810
rect 27234 3189 32856 3190
rect 26944 3062 27071 3078
rect 32963 3078 33010 8922
rect 33074 3078 33090 8922
rect 38982 8922 39109 8938
rect 33253 8810 38875 8811
rect 33253 3190 33254 8810
rect 38874 3190 38875 8810
rect 33253 3189 38875 3190
rect 32963 3062 33090 3078
rect 38982 3078 39029 8922
rect 39093 3078 39109 8922
rect 45001 8922 45128 8938
rect 39272 8810 44894 8811
rect 39272 3190 39273 8810
rect 44893 3190 44894 8810
rect 39272 3189 44894 3190
rect 38982 3062 39109 3078
rect 45001 3078 45048 8922
rect 45112 3078 45128 8922
rect 45001 3062 45128 3078
rect -39265 2938 -39161 3062
rect -33246 2938 -33142 3062
rect -27227 2938 -27123 3062
rect -21208 2938 -21104 3062
rect -15189 2938 -15085 3062
rect -9170 2938 -9066 3062
rect -3151 2938 -3047 3062
rect 2868 2938 2972 3062
rect 8887 2938 8991 3062
rect 14906 2938 15010 3062
rect 20925 2938 21029 3062
rect 26944 2938 27048 3062
rect 32963 2938 33067 3062
rect 38982 2938 39086 3062
rect 45001 2938 45105 3062
rect -39265 2922 -39138 2938
rect -44994 2810 -39372 2811
rect -44994 -2810 -44993 2810
rect -39373 -2810 -39372 2810
rect -44994 -2811 -39372 -2810
rect -39265 -2922 -39218 2922
rect -39154 -2922 -39138 2922
rect -33246 2922 -33119 2938
rect -38975 2810 -33353 2811
rect -38975 -2810 -38974 2810
rect -33354 -2810 -33353 2810
rect -38975 -2811 -33353 -2810
rect -39265 -2938 -39138 -2922
rect -33246 -2922 -33199 2922
rect -33135 -2922 -33119 2922
rect -27227 2922 -27100 2938
rect -32956 2810 -27334 2811
rect -32956 -2810 -32955 2810
rect -27335 -2810 -27334 2810
rect -32956 -2811 -27334 -2810
rect -33246 -2938 -33119 -2922
rect -27227 -2922 -27180 2922
rect -27116 -2922 -27100 2922
rect -21208 2922 -21081 2938
rect -26937 2810 -21315 2811
rect -26937 -2810 -26936 2810
rect -21316 -2810 -21315 2810
rect -26937 -2811 -21315 -2810
rect -27227 -2938 -27100 -2922
rect -21208 -2922 -21161 2922
rect -21097 -2922 -21081 2922
rect -15189 2922 -15062 2938
rect -20918 2810 -15296 2811
rect -20918 -2810 -20917 2810
rect -15297 -2810 -15296 2810
rect -20918 -2811 -15296 -2810
rect -21208 -2938 -21081 -2922
rect -15189 -2922 -15142 2922
rect -15078 -2922 -15062 2922
rect -9170 2922 -9043 2938
rect -14899 2810 -9277 2811
rect -14899 -2810 -14898 2810
rect -9278 -2810 -9277 2810
rect -14899 -2811 -9277 -2810
rect -15189 -2938 -15062 -2922
rect -9170 -2922 -9123 2922
rect -9059 -2922 -9043 2922
rect -3151 2922 -3024 2938
rect -8880 2810 -3258 2811
rect -8880 -2810 -8879 2810
rect -3259 -2810 -3258 2810
rect -8880 -2811 -3258 -2810
rect -9170 -2938 -9043 -2922
rect -3151 -2922 -3104 2922
rect -3040 -2922 -3024 2922
rect 2868 2922 2995 2938
rect -2861 2810 2761 2811
rect -2861 -2810 -2860 2810
rect 2760 -2810 2761 2810
rect -2861 -2811 2761 -2810
rect -3151 -2938 -3024 -2922
rect 2868 -2922 2915 2922
rect 2979 -2922 2995 2922
rect 8887 2922 9014 2938
rect 3158 2810 8780 2811
rect 3158 -2810 3159 2810
rect 8779 -2810 8780 2810
rect 3158 -2811 8780 -2810
rect 2868 -2938 2995 -2922
rect 8887 -2922 8934 2922
rect 8998 -2922 9014 2922
rect 14906 2922 15033 2938
rect 9177 2810 14799 2811
rect 9177 -2810 9178 2810
rect 14798 -2810 14799 2810
rect 9177 -2811 14799 -2810
rect 8887 -2938 9014 -2922
rect 14906 -2922 14953 2922
rect 15017 -2922 15033 2922
rect 20925 2922 21052 2938
rect 15196 2810 20818 2811
rect 15196 -2810 15197 2810
rect 20817 -2810 20818 2810
rect 15196 -2811 20818 -2810
rect 14906 -2938 15033 -2922
rect 20925 -2922 20972 2922
rect 21036 -2922 21052 2922
rect 26944 2922 27071 2938
rect 21215 2810 26837 2811
rect 21215 -2810 21216 2810
rect 26836 -2810 26837 2810
rect 21215 -2811 26837 -2810
rect 20925 -2938 21052 -2922
rect 26944 -2922 26991 2922
rect 27055 -2922 27071 2922
rect 32963 2922 33090 2938
rect 27234 2810 32856 2811
rect 27234 -2810 27235 2810
rect 32855 -2810 32856 2810
rect 27234 -2811 32856 -2810
rect 26944 -2938 27071 -2922
rect 32963 -2922 33010 2922
rect 33074 -2922 33090 2922
rect 38982 2922 39109 2938
rect 33253 2810 38875 2811
rect 33253 -2810 33254 2810
rect 38874 -2810 38875 2810
rect 33253 -2811 38875 -2810
rect 32963 -2938 33090 -2922
rect 38982 -2922 39029 2922
rect 39093 -2922 39109 2922
rect 45001 2922 45128 2938
rect 39272 2810 44894 2811
rect 39272 -2810 39273 2810
rect 44893 -2810 44894 2810
rect 39272 -2811 44894 -2810
rect 38982 -2938 39109 -2922
rect 45001 -2922 45048 2922
rect 45112 -2922 45128 2922
rect 45001 -2938 45128 -2922
rect -39265 -3062 -39161 -2938
rect -33246 -3062 -33142 -2938
rect -27227 -3062 -27123 -2938
rect -21208 -3062 -21104 -2938
rect -15189 -3062 -15085 -2938
rect -9170 -3062 -9066 -2938
rect -3151 -3062 -3047 -2938
rect 2868 -3062 2972 -2938
rect 8887 -3062 8991 -2938
rect 14906 -3062 15010 -2938
rect 20925 -3062 21029 -2938
rect 26944 -3062 27048 -2938
rect 32963 -3062 33067 -2938
rect 38982 -3062 39086 -2938
rect 45001 -3062 45105 -2938
rect -39265 -3078 -39138 -3062
rect -44994 -3190 -39372 -3189
rect -44994 -8810 -44993 -3190
rect -39373 -8810 -39372 -3190
rect -44994 -8811 -39372 -8810
rect -39265 -8922 -39218 -3078
rect -39154 -8922 -39138 -3078
rect -33246 -3078 -33119 -3062
rect -38975 -3190 -33353 -3189
rect -38975 -8810 -38974 -3190
rect -33354 -8810 -33353 -3190
rect -38975 -8811 -33353 -8810
rect -39265 -8938 -39138 -8922
rect -33246 -8922 -33199 -3078
rect -33135 -8922 -33119 -3078
rect -27227 -3078 -27100 -3062
rect -32956 -3190 -27334 -3189
rect -32956 -8810 -32955 -3190
rect -27335 -8810 -27334 -3190
rect -32956 -8811 -27334 -8810
rect -33246 -8938 -33119 -8922
rect -27227 -8922 -27180 -3078
rect -27116 -8922 -27100 -3078
rect -21208 -3078 -21081 -3062
rect -26937 -3190 -21315 -3189
rect -26937 -8810 -26936 -3190
rect -21316 -8810 -21315 -3190
rect -26937 -8811 -21315 -8810
rect -27227 -8938 -27100 -8922
rect -21208 -8922 -21161 -3078
rect -21097 -8922 -21081 -3078
rect -15189 -3078 -15062 -3062
rect -20918 -3190 -15296 -3189
rect -20918 -8810 -20917 -3190
rect -15297 -8810 -15296 -3190
rect -20918 -8811 -15296 -8810
rect -21208 -8938 -21081 -8922
rect -15189 -8922 -15142 -3078
rect -15078 -8922 -15062 -3078
rect -9170 -3078 -9043 -3062
rect -14899 -3190 -9277 -3189
rect -14899 -8810 -14898 -3190
rect -9278 -8810 -9277 -3190
rect -14899 -8811 -9277 -8810
rect -15189 -8938 -15062 -8922
rect -9170 -8922 -9123 -3078
rect -9059 -8922 -9043 -3078
rect -3151 -3078 -3024 -3062
rect -8880 -3190 -3258 -3189
rect -8880 -8810 -8879 -3190
rect -3259 -8810 -3258 -3190
rect -8880 -8811 -3258 -8810
rect -9170 -8938 -9043 -8922
rect -3151 -8922 -3104 -3078
rect -3040 -8922 -3024 -3078
rect 2868 -3078 2995 -3062
rect -2861 -3190 2761 -3189
rect -2861 -8810 -2860 -3190
rect 2760 -8810 2761 -3190
rect -2861 -8811 2761 -8810
rect -3151 -8938 -3024 -8922
rect 2868 -8922 2915 -3078
rect 2979 -8922 2995 -3078
rect 8887 -3078 9014 -3062
rect 3158 -3190 8780 -3189
rect 3158 -8810 3159 -3190
rect 8779 -8810 8780 -3190
rect 3158 -8811 8780 -8810
rect 2868 -8938 2995 -8922
rect 8887 -8922 8934 -3078
rect 8998 -8922 9014 -3078
rect 14906 -3078 15033 -3062
rect 9177 -3190 14799 -3189
rect 9177 -8810 9178 -3190
rect 14798 -8810 14799 -3190
rect 9177 -8811 14799 -8810
rect 8887 -8938 9014 -8922
rect 14906 -8922 14953 -3078
rect 15017 -8922 15033 -3078
rect 20925 -3078 21052 -3062
rect 15196 -3190 20818 -3189
rect 15196 -8810 15197 -3190
rect 20817 -8810 20818 -3190
rect 15196 -8811 20818 -8810
rect 14906 -8938 15033 -8922
rect 20925 -8922 20972 -3078
rect 21036 -8922 21052 -3078
rect 26944 -3078 27071 -3062
rect 21215 -3190 26837 -3189
rect 21215 -8810 21216 -3190
rect 26836 -8810 26837 -3190
rect 21215 -8811 26837 -8810
rect 20925 -8938 21052 -8922
rect 26944 -8922 26991 -3078
rect 27055 -8922 27071 -3078
rect 32963 -3078 33090 -3062
rect 27234 -3190 32856 -3189
rect 27234 -8810 27235 -3190
rect 32855 -8810 32856 -3190
rect 27234 -8811 32856 -8810
rect 26944 -8938 27071 -8922
rect 32963 -8922 33010 -3078
rect 33074 -8922 33090 -3078
rect 38982 -3078 39109 -3062
rect 33253 -3190 38875 -3189
rect 33253 -8810 33254 -3190
rect 38874 -8810 38875 -3190
rect 33253 -8811 38875 -8810
rect 32963 -8938 33090 -8922
rect 38982 -8922 39029 -3078
rect 39093 -8922 39109 -3078
rect 45001 -3078 45128 -3062
rect 39272 -3190 44894 -3189
rect 39272 -8810 39273 -3190
rect 44893 -8810 44894 -3190
rect 39272 -8811 44894 -8810
rect 38982 -8938 39109 -8922
rect 45001 -8922 45048 -3078
rect 45112 -8922 45128 -3078
rect 45001 -8938 45128 -8922
rect -39265 -9062 -39161 -8938
rect -33246 -9062 -33142 -8938
rect -27227 -9062 -27123 -8938
rect -21208 -9062 -21104 -8938
rect -15189 -9062 -15085 -8938
rect -9170 -9062 -9066 -8938
rect -3151 -9062 -3047 -8938
rect 2868 -9062 2972 -8938
rect 8887 -9062 8991 -8938
rect 14906 -9062 15010 -8938
rect 20925 -9062 21029 -8938
rect 26944 -9062 27048 -8938
rect 32963 -9062 33067 -8938
rect 38982 -9062 39086 -8938
rect 45001 -9062 45105 -8938
rect -39265 -9078 -39138 -9062
rect -44994 -9190 -39372 -9189
rect -44994 -14810 -44993 -9190
rect -39373 -14810 -39372 -9190
rect -44994 -14811 -39372 -14810
rect -39265 -14922 -39218 -9078
rect -39154 -14922 -39138 -9078
rect -33246 -9078 -33119 -9062
rect -38975 -9190 -33353 -9189
rect -38975 -14810 -38974 -9190
rect -33354 -14810 -33353 -9190
rect -38975 -14811 -33353 -14810
rect -39265 -14938 -39138 -14922
rect -33246 -14922 -33199 -9078
rect -33135 -14922 -33119 -9078
rect -27227 -9078 -27100 -9062
rect -32956 -9190 -27334 -9189
rect -32956 -14810 -32955 -9190
rect -27335 -14810 -27334 -9190
rect -32956 -14811 -27334 -14810
rect -33246 -14938 -33119 -14922
rect -27227 -14922 -27180 -9078
rect -27116 -14922 -27100 -9078
rect -21208 -9078 -21081 -9062
rect -26937 -9190 -21315 -9189
rect -26937 -14810 -26936 -9190
rect -21316 -14810 -21315 -9190
rect -26937 -14811 -21315 -14810
rect -27227 -14938 -27100 -14922
rect -21208 -14922 -21161 -9078
rect -21097 -14922 -21081 -9078
rect -15189 -9078 -15062 -9062
rect -20918 -9190 -15296 -9189
rect -20918 -14810 -20917 -9190
rect -15297 -14810 -15296 -9190
rect -20918 -14811 -15296 -14810
rect -21208 -14938 -21081 -14922
rect -15189 -14922 -15142 -9078
rect -15078 -14922 -15062 -9078
rect -9170 -9078 -9043 -9062
rect -14899 -9190 -9277 -9189
rect -14899 -14810 -14898 -9190
rect -9278 -14810 -9277 -9190
rect -14899 -14811 -9277 -14810
rect -15189 -14938 -15062 -14922
rect -9170 -14922 -9123 -9078
rect -9059 -14922 -9043 -9078
rect -3151 -9078 -3024 -9062
rect -8880 -9190 -3258 -9189
rect -8880 -14810 -8879 -9190
rect -3259 -14810 -3258 -9190
rect -8880 -14811 -3258 -14810
rect -9170 -14938 -9043 -14922
rect -3151 -14922 -3104 -9078
rect -3040 -14922 -3024 -9078
rect 2868 -9078 2995 -9062
rect -2861 -9190 2761 -9189
rect -2861 -14810 -2860 -9190
rect 2760 -14810 2761 -9190
rect -2861 -14811 2761 -14810
rect -3151 -14938 -3024 -14922
rect 2868 -14922 2915 -9078
rect 2979 -14922 2995 -9078
rect 8887 -9078 9014 -9062
rect 3158 -9190 8780 -9189
rect 3158 -14810 3159 -9190
rect 8779 -14810 8780 -9190
rect 3158 -14811 8780 -14810
rect 2868 -14938 2995 -14922
rect 8887 -14922 8934 -9078
rect 8998 -14922 9014 -9078
rect 14906 -9078 15033 -9062
rect 9177 -9190 14799 -9189
rect 9177 -14810 9178 -9190
rect 14798 -14810 14799 -9190
rect 9177 -14811 14799 -14810
rect 8887 -14938 9014 -14922
rect 14906 -14922 14953 -9078
rect 15017 -14922 15033 -9078
rect 20925 -9078 21052 -9062
rect 15196 -9190 20818 -9189
rect 15196 -14810 15197 -9190
rect 20817 -14810 20818 -9190
rect 15196 -14811 20818 -14810
rect 14906 -14938 15033 -14922
rect 20925 -14922 20972 -9078
rect 21036 -14922 21052 -9078
rect 26944 -9078 27071 -9062
rect 21215 -9190 26837 -9189
rect 21215 -14810 21216 -9190
rect 26836 -14810 26837 -9190
rect 21215 -14811 26837 -14810
rect 20925 -14938 21052 -14922
rect 26944 -14922 26991 -9078
rect 27055 -14922 27071 -9078
rect 32963 -9078 33090 -9062
rect 27234 -9190 32856 -9189
rect 27234 -14810 27235 -9190
rect 32855 -14810 32856 -9190
rect 27234 -14811 32856 -14810
rect 26944 -14938 27071 -14922
rect 32963 -14922 33010 -9078
rect 33074 -14922 33090 -9078
rect 38982 -9078 39109 -9062
rect 33253 -9190 38875 -9189
rect 33253 -14810 33254 -9190
rect 38874 -14810 38875 -9190
rect 33253 -14811 38875 -14810
rect 32963 -14938 33090 -14922
rect 38982 -14922 39029 -9078
rect 39093 -14922 39109 -9078
rect 45001 -9078 45128 -9062
rect 39272 -9190 44894 -9189
rect 39272 -14810 39273 -9190
rect 44893 -14810 44894 -9190
rect 39272 -14811 44894 -14810
rect 38982 -14938 39109 -14922
rect 45001 -14922 45048 -9078
rect 45112 -14922 45128 -9078
rect 45001 -14938 45128 -14922
rect -39265 -15062 -39161 -14938
rect -33246 -15062 -33142 -14938
rect -27227 -15062 -27123 -14938
rect -21208 -15062 -21104 -14938
rect -15189 -15062 -15085 -14938
rect -9170 -15062 -9066 -14938
rect -3151 -15062 -3047 -14938
rect 2868 -15062 2972 -14938
rect 8887 -15062 8991 -14938
rect 14906 -15062 15010 -14938
rect 20925 -15062 21029 -14938
rect 26944 -15062 27048 -14938
rect 32963 -15062 33067 -14938
rect 38982 -15062 39086 -14938
rect 45001 -15062 45105 -14938
rect -39265 -15078 -39138 -15062
rect -44994 -15190 -39372 -15189
rect -44994 -20810 -44993 -15190
rect -39373 -20810 -39372 -15190
rect -44994 -20811 -39372 -20810
rect -39265 -20922 -39218 -15078
rect -39154 -20922 -39138 -15078
rect -33246 -15078 -33119 -15062
rect -38975 -15190 -33353 -15189
rect -38975 -20810 -38974 -15190
rect -33354 -20810 -33353 -15190
rect -38975 -20811 -33353 -20810
rect -39265 -20938 -39138 -20922
rect -33246 -20922 -33199 -15078
rect -33135 -20922 -33119 -15078
rect -27227 -15078 -27100 -15062
rect -32956 -15190 -27334 -15189
rect -32956 -20810 -32955 -15190
rect -27335 -20810 -27334 -15190
rect -32956 -20811 -27334 -20810
rect -33246 -20938 -33119 -20922
rect -27227 -20922 -27180 -15078
rect -27116 -20922 -27100 -15078
rect -21208 -15078 -21081 -15062
rect -26937 -15190 -21315 -15189
rect -26937 -20810 -26936 -15190
rect -21316 -20810 -21315 -15190
rect -26937 -20811 -21315 -20810
rect -27227 -20938 -27100 -20922
rect -21208 -20922 -21161 -15078
rect -21097 -20922 -21081 -15078
rect -15189 -15078 -15062 -15062
rect -20918 -15190 -15296 -15189
rect -20918 -20810 -20917 -15190
rect -15297 -20810 -15296 -15190
rect -20918 -20811 -15296 -20810
rect -21208 -20938 -21081 -20922
rect -15189 -20922 -15142 -15078
rect -15078 -20922 -15062 -15078
rect -9170 -15078 -9043 -15062
rect -14899 -15190 -9277 -15189
rect -14899 -20810 -14898 -15190
rect -9278 -20810 -9277 -15190
rect -14899 -20811 -9277 -20810
rect -15189 -20938 -15062 -20922
rect -9170 -20922 -9123 -15078
rect -9059 -20922 -9043 -15078
rect -3151 -15078 -3024 -15062
rect -8880 -15190 -3258 -15189
rect -8880 -20810 -8879 -15190
rect -3259 -20810 -3258 -15190
rect -8880 -20811 -3258 -20810
rect -9170 -20938 -9043 -20922
rect -3151 -20922 -3104 -15078
rect -3040 -20922 -3024 -15078
rect 2868 -15078 2995 -15062
rect -2861 -15190 2761 -15189
rect -2861 -20810 -2860 -15190
rect 2760 -20810 2761 -15190
rect -2861 -20811 2761 -20810
rect -3151 -20938 -3024 -20922
rect 2868 -20922 2915 -15078
rect 2979 -20922 2995 -15078
rect 8887 -15078 9014 -15062
rect 3158 -15190 8780 -15189
rect 3158 -20810 3159 -15190
rect 8779 -20810 8780 -15190
rect 3158 -20811 8780 -20810
rect 2868 -20938 2995 -20922
rect 8887 -20922 8934 -15078
rect 8998 -20922 9014 -15078
rect 14906 -15078 15033 -15062
rect 9177 -15190 14799 -15189
rect 9177 -20810 9178 -15190
rect 14798 -20810 14799 -15190
rect 9177 -20811 14799 -20810
rect 8887 -20938 9014 -20922
rect 14906 -20922 14953 -15078
rect 15017 -20922 15033 -15078
rect 20925 -15078 21052 -15062
rect 15196 -15190 20818 -15189
rect 15196 -20810 15197 -15190
rect 20817 -20810 20818 -15190
rect 15196 -20811 20818 -20810
rect 14906 -20938 15033 -20922
rect 20925 -20922 20972 -15078
rect 21036 -20922 21052 -15078
rect 26944 -15078 27071 -15062
rect 21215 -15190 26837 -15189
rect 21215 -20810 21216 -15190
rect 26836 -20810 26837 -15190
rect 21215 -20811 26837 -20810
rect 20925 -20938 21052 -20922
rect 26944 -20922 26991 -15078
rect 27055 -20922 27071 -15078
rect 32963 -15078 33090 -15062
rect 27234 -15190 32856 -15189
rect 27234 -20810 27235 -15190
rect 32855 -20810 32856 -15190
rect 27234 -20811 32856 -20810
rect 26944 -20938 27071 -20922
rect 32963 -20922 33010 -15078
rect 33074 -20922 33090 -15078
rect 38982 -15078 39109 -15062
rect 33253 -15190 38875 -15189
rect 33253 -20810 33254 -15190
rect 38874 -20810 38875 -15190
rect 33253 -20811 38875 -20810
rect 32963 -20938 33090 -20922
rect 38982 -20922 39029 -15078
rect 39093 -20922 39109 -15078
rect 45001 -15078 45128 -15062
rect 39272 -15190 44894 -15189
rect 39272 -20810 39273 -15190
rect 44893 -20810 44894 -15190
rect 39272 -20811 44894 -20810
rect 38982 -20938 39109 -20922
rect 45001 -20922 45048 -15078
rect 45112 -20922 45128 -15078
rect 45001 -20938 45128 -20922
rect -39265 -21000 -39161 -20938
rect -33246 -21000 -33142 -20938
rect -27227 -21000 -27123 -20938
rect -21208 -21000 -21104 -20938
rect -15189 -21000 -15085 -20938
rect -9170 -21000 -9066 -20938
rect -3151 -21000 -3047 -20938
rect 2868 -21000 2972 -20938
rect 8887 -21000 8991 -20938
rect 14906 -21000 15010 -20938
rect 20925 -21000 21029 -20938
rect 26944 -21000 27048 -20938
rect 32963 -21000 33067 -20938
rect 38982 -21000 39086 -20938
rect 45001 -21000 45105 -20938
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX 39133 15050 45033 20950
string parameters w 28.5 l 28.5 val 1.646k carea 2.00 cperi 0.19 nx 15 ny 7 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 0 ccov 100
string library sky130
<< end >>
