magic
tech sky130A
magscale 1 2
timestamp 1634373541
<< pwell >>
rect 36 -10642 388 -10336
rect 226 -19826 392 -19276
rect -582 -20056 682 -19826
rect 46 -20498 454 -20246
<< locali >>
rect 430 9308 504 9334
rect 430 9250 438 9308
rect 494 9250 504 9308
rect 430 9202 504 9250
rect 496 -298 574 -282
rect 496 -376 504 -298
rect 566 -376 574 -298
rect 496 -396 574 -376
rect 16304 -10082 16428 -10040
rect 16304 -10186 16322 -10082
rect 16408 -10186 16428 -10082
rect 16304 -10212 16428 -10186
rect 16268 -19898 16496 -19756
rect 16268 -20086 16320 -19898
rect 16450 -20086 16496 -19898
rect 16268 -20106 16496 -20086
<< viali >>
rect 438 9250 494 9308
rect 504 -376 566 -298
rect 16322 -10186 16408 -10082
rect 16320 -20086 16450 -19898
<< metal1 >>
rect 16366 9344 16582 9474
rect 432 9308 504 9334
rect 432 9250 438 9308
rect 494 9250 504 9308
rect 432 9238 504 9250
rect -14 -166 198 354
rect -14 -238 20 -166
rect 172 -238 198 -166
rect -14 -248 198 -238
rect 290 144 432 174
rect 290 12 508 144
rect 290 -76 514 12
rect -910 -1034 210 -482
rect 290 -504 432 -76
rect 496 -298 574 -282
rect 496 -376 504 -298
rect 566 -376 574 -298
rect 496 -396 574 -376
rect 74 -9936 272 -9304
rect 74 -10056 606 -9936
rect 16304 -10082 16428 -10040
rect 532 -10216 556 -10130
rect 16304 -10186 16322 -10082
rect 16408 -10186 16428 -10082
rect 16304 -10212 16428 -10186
rect 36 -10416 388 -10336
rect 36 -10572 74 -10416
rect 198 -10572 388 -10416
rect 36 -10642 388 -10572
rect 226 -19826 392 -19276
rect -582 -19862 682 -19826
rect -582 -20030 -564 -19862
rect -378 -20030 682 -19862
rect -582 -20056 682 -20030
rect 16268 -19898 16496 -19756
rect 16268 -20086 16320 -19898
rect 16450 -20086 16496 -19898
rect 16268 -20106 16496 -20086
rect 46 -20292 454 -20246
rect 46 -20476 68 -20292
rect 194 -20476 454 -20292
rect 46 -20498 454 -20476
<< via1 >>
rect 438 9250 494 9308
rect 20 -238 172 -166
rect 504 -376 566 -298
rect 16322 -10186 16408 -10082
rect 74 -10572 198 -10416
rect -564 -20030 -378 -19862
rect 16320 -20086 16450 -19898
rect 68 -20476 194 -20292
<< metal2 >>
rect -654 -114 -342 -110
rect -724 -144 224 -114
rect -724 -166 580 -144
rect -724 -238 20 -166
rect 172 -238 580 -166
rect -724 -248 580 -238
rect -724 -316 224 -248
rect -654 -19862 -342 -316
rect 16370 -446 16498 440
rect 404 -9654 662 -9382
rect -40 -9664 672 -9654
rect -42 -9862 672 -9664
rect -42 -9908 202 -9862
rect -42 -10416 214 -9908
rect 16292 -10082 17472 -9840
rect 16292 -10156 16322 -10082
rect 16408 -10156 17472 -10082
rect -42 -10444 74 -10416
rect -30 -10572 74 -10444
rect 198 -10450 214 -10416
rect 198 -10572 398 -10450
rect -30 -10688 398 -10572
rect 416 -19582 580 -18916
rect -654 -20030 -564 -19862
rect -378 -20030 -342 -19862
rect -654 -20060 -342 -20030
rect 32 -19770 590 -19582
rect 16270 -19754 16492 -19226
rect 32 -20292 232 -19770
rect 16270 -19898 16496 -19754
rect 16270 -20024 16320 -19898
rect 16276 -20086 16320 -20024
rect 16450 -20086 16496 -19898
rect 16276 -20112 16496 -20086
rect 32 -20476 68 -20292
rect 194 -20476 232 -20292
rect 32 -20498 232 -20476
use pmos20  pmos20_0
timestamp 1634295700
transform 0 1 266 -1 0 9220
box -238 -278 9216 16385
use pmos20  pmos20_1
timestamp 1634295700
transform 0 1 334 -1 0 -342
box -238 -278 9216 16385
use nmos20  nmos20_1
timestamp 1634288453
transform 0 -1 8575 -1 0 -20124
box -308 -8222 9194 8295
use nmos20  nmos20_0
timestamp 1634288453
transform 0 -1 8511 -1 0 -10210
box -308 -8222 9194 8295
<< labels >>
rlabel metal1 16536 9384 16536 9384 1 VIN1
rlabel metal2 17042 -10074 17042 -10074 1 VSS
rlabel via1 -426 -19954 -426 -19954 1 VINN
rlabel metal1 -146 -846 -146 -846 1 VINP
<< end >>
