magic
tech sky130A
magscale 1 2
timestamp 1634206901
<< error_p >>
rect -31 5081 31 5087
rect -31 5047 -19 5081
rect -31 5041 31 5047
rect -31 -5047 31 -5041
rect -31 -5081 -19 -5047
rect -31 -5087 31 -5081
<< nwell >>
rect -231 -5219 231 5219
<< pmoslvt >>
rect -35 -5000 35 5000
<< pdiff >>
rect -93 4988 -35 5000
rect -93 -4988 -81 4988
rect -47 -4988 -35 4988
rect -93 -5000 -35 -4988
rect 35 4988 93 5000
rect 35 -4988 47 4988
rect 81 -4988 93 4988
rect 35 -5000 93 -4988
<< pdiffc >>
rect -81 -4988 -47 4988
rect 47 -4988 81 4988
<< nsubdiff >>
rect -195 5149 -99 5183
rect 99 5149 195 5183
rect -195 5087 -161 5149
rect 161 5087 195 5149
rect -195 -5149 -161 -5087
rect 161 -5149 195 -5087
rect -195 -5183 -99 -5149
rect 99 -5183 195 -5149
<< nsubdiffcont >>
rect -99 5149 99 5183
rect -195 -5087 -161 5087
rect 161 -5087 195 5087
rect -99 -5183 99 -5149
<< poly >>
rect -35 5081 35 5097
rect -35 5047 -19 5081
rect 19 5047 35 5081
rect -35 5000 35 5047
rect -35 -5047 35 -5000
rect -35 -5081 -19 -5047
rect 19 -5081 35 -5047
rect -35 -5097 35 -5081
<< polycont >>
rect -19 5047 19 5081
rect -19 -5081 19 -5047
<< locali >>
rect -195 5149 -99 5183
rect 99 5149 195 5183
rect -195 5087 -161 5149
rect 161 5087 195 5149
rect -35 5047 -19 5081
rect 19 5047 35 5081
rect -81 4988 -47 5004
rect -81 -5004 -47 -4988
rect 47 4988 81 5004
rect 47 -5004 81 -4988
rect -35 -5081 -19 -5047
rect 19 -5081 35 -5047
rect -195 -5149 -161 -5087
rect 161 -5149 195 -5087
rect -195 -5183 -99 -5149
rect 99 -5183 195 -5149
<< viali >>
rect -19 5047 19 5081
rect -81 -4988 -47 4988
rect 47 -4988 81 4988
rect -19 -5081 19 -5047
<< metal1 >>
rect -31 5081 31 5087
rect -31 5047 -19 5081
rect 19 5047 31 5081
rect -31 5041 31 5047
rect -87 4988 -41 5000
rect -87 -4988 -81 4988
rect -47 -4988 -41 4988
rect -87 -5000 -41 -4988
rect 41 4988 87 5000
rect 41 -4988 47 4988
rect 81 -4988 87 4988
rect 41 -5000 87 -4988
rect -31 -5047 31 -5041
rect -31 -5081 -19 -5047
rect 19 -5081 31 -5047
rect -31 -5087 31 -5081
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string FIXED_BBOX -178 -5166 178 5166
string parameters w 50 l 0.35 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
