magic
tech sky130A
magscale 1 2
timestamp 1634294201
<< error_p >>
rect -41144 41000 -41084 47200
rect -41064 41000 -41004 47200
rect -34825 41000 -34765 47200
rect -34745 41000 -34685 47200
rect -28506 41000 -28446 47200
rect -28426 41000 -28366 47200
rect -22187 41000 -22127 47200
rect -22107 41000 -22047 47200
rect -15868 41000 -15808 47200
rect -15788 41000 -15728 47200
rect -9549 41000 -9489 47200
rect -9469 41000 -9409 47200
rect -3230 41000 -3170 47200
rect -3150 41000 -3090 47200
rect 3089 41000 3149 47200
rect 3169 41000 3229 47200
rect 9408 41000 9468 47200
rect 9488 41000 9548 47200
rect 15727 41000 15787 47200
rect 15807 41000 15867 47200
rect 22046 41000 22106 47200
rect 22126 41000 22186 47200
rect 28365 41000 28425 47200
rect 28445 41000 28505 47200
rect 34684 41000 34744 47200
rect 34764 41000 34824 47200
rect 41003 41000 41063 47200
rect 41083 41000 41143 47200
rect -41144 34700 -41084 40900
rect -41064 34700 -41004 40900
rect -34825 34700 -34765 40900
rect -34745 34700 -34685 40900
rect -28506 34700 -28446 40900
rect -28426 34700 -28366 40900
rect -22187 34700 -22127 40900
rect -22107 34700 -22047 40900
rect -15868 34700 -15808 40900
rect -15788 34700 -15728 40900
rect -9549 34700 -9489 40900
rect -9469 34700 -9409 40900
rect -3230 34700 -3170 40900
rect -3150 34700 -3090 40900
rect 3089 34700 3149 40900
rect 3169 34700 3229 40900
rect 9408 34700 9468 40900
rect 9488 34700 9548 40900
rect 15727 34700 15787 40900
rect 15807 34700 15867 40900
rect 22046 34700 22106 40900
rect 22126 34700 22186 40900
rect 28365 34700 28425 40900
rect 28445 34700 28505 40900
rect 34684 34700 34744 40900
rect 34764 34700 34824 40900
rect 41003 34700 41063 40900
rect 41083 34700 41143 40900
rect -41144 28400 -41084 34600
rect -41064 28400 -41004 34600
rect -34825 28400 -34765 34600
rect -34745 28400 -34685 34600
rect -28506 28400 -28446 34600
rect -28426 28400 -28366 34600
rect -22187 28400 -22127 34600
rect -22107 28400 -22047 34600
rect -15868 28400 -15808 34600
rect -15788 28400 -15728 34600
rect -9549 28400 -9489 34600
rect -9469 28400 -9409 34600
rect -3230 28400 -3170 34600
rect -3150 28400 -3090 34600
rect 3089 28400 3149 34600
rect 3169 28400 3229 34600
rect 9408 28400 9468 34600
rect 9488 28400 9548 34600
rect 15727 28400 15787 34600
rect 15807 28400 15867 34600
rect 22046 28400 22106 34600
rect 22126 28400 22186 34600
rect 28365 28400 28425 34600
rect 28445 28400 28505 34600
rect 34684 28400 34744 34600
rect 34764 28400 34824 34600
rect 41003 28400 41063 34600
rect 41083 28400 41143 34600
rect -41144 22100 -41084 28300
rect -41064 22100 -41004 28300
rect -34825 22100 -34765 28300
rect -34745 22100 -34685 28300
rect -28506 22100 -28446 28300
rect -28426 22100 -28366 28300
rect -22187 22100 -22127 28300
rect -22107 22100 -22047 28300
rect -15868 22100 -15808 28300
rect -15788 22100 -15728 28300
rect -9549 22100 -9489 28300
rect -9469 22100 -9409 28300
rect -3230 22100 -3170 28300
rect -3150 22100 -3090 28300
rect 3089 22100 3149 28300
rect 3169 22100 3229 28300
rect 9408 22100 9468 28300
rect 9488 22100 9548 28300
rect 15727 22100 15787 28300
rect 15807 22100 15867 28300
rect 22046 22100 22106 28300
rect 22126 22100 22186 28300
rect 28365 22100 28425 28300
rect 28445 22100 28505 28300
rect 34684 22100 34744 28300
rect 34764 22100 34824 28300
rect 41003 22100 41063 28300
rect 41083 22100 41143 28300
rect -41144 15800 -41084 22000
rect -41064 15800 -41004 22000
rect -34825 15800 -34765 22000
rect -34745 15800 -34685 22000
rect -28506 15800 -28446 22000
rect -28426 15800 -28366 22000
rect -22187 15800 -22127 22000
rect -22107 15800 -22047 22000
rect -15868 15800 -15808 22000
rect -15788 15800 -15728 22000
rect -9549 15800 -9489 22000
rect -9469 15800 -9409 22000
rect -3230 15800 -3170 22000
rect -3150 15800 -3090 22000
rect 3089 15800 3149 22000
rect 3169 15800 3229 22000
rect 9408 15800 9468 22000
rect 9488 15800 9548 22000
rect 15727 15800 15787 22000
rect 15807 15800 15867 22000
rect 22046 15800 22106 22000
rect 22126 15800 22186 22000
rect 28365 15800 28425 22000
rect 28445 15800 28505 22000
rect 34684 15800 34744 22000
rect 34764 15800 34824 22000
rect 41003 15800 41063 22000
rect 41083 15800 41143 22000
rect -41144 9500 -41084 15700
rect -41064 9500 -41004 15700
rect -34825 9500 -34765 15700
rect -34745 9500 -34685 15700
rect -28506 9500 -28446 15700
rect -28426 9500 -28366 15700
rect -22187 9500 -22127 15700
rect -22107 9500 -22047 15700
rect -15868 9500 -15808 15700
rect -15788 9500 -15728 15700
rect -9549 9500 -9489 15700
rect -9469 9500 -9409 15700
rect -3230 9500 -3170 15700
rect -3150 9500 -3090 15700
rect 3089 9500 3149 15700
rect 3169 9500 3229 15700
rect 9408 9500 9468 15700
rect 9488 9500 9548 15700
rect 15727 9500 15787 15700
rect 15807 9500 15867 15700
rect 22046 9500 22106 15700
rect 22126 9500 22186 15700
rect 28365 9500 28425 15700
rect 28445 9500 28505 15700
rect 34684 9500 34744 15700
rect 34764 9500 34824 15700
rect 41003 9500 41063 15700
rect 41083 9500 41143 15700
rect -41144 3200 -41084 9400
rect -41064 3200 -41004 9400
rect -34825 3200 -34765 9400
rect -34745 3200 -34685 9400
rect -28506 3200 -28446 9400
rect -28426 3200 -28366 9400
rect -22187 3200 -22127 9400
rect -22107 3200 -22047 9400
rect -15868 3200 -15808 9400
rect -15788 3200 -15728 9400
rect -9549 3200 -9489 9400
rect -9469 3200 -9409 9400
rect -3230 3200 -3170 9400
rect -3150 3200 -3090 9400
rect 3089 3200 3149 9400
rect 3169 3200 3229 9400
rect 9408 3200 9468 9400
rect 9488 3200 9548 9400
rect 15727 3200 15787 9400
rect 15807 3200 15867 9400
rect 22046 3200 22106 9400
rect 22126 3200 22186 9400
rect 28365 3200 28425 9400
rect 28445 3200 28505 9400
rect 34684 3200 34744 9400
rect 34764 3200 34824 9400
rect 41003 3200 41063 9400
rect 41083 3200 41143 9400
rect -41144 -3100 -41084 3100
rect -41064 -3100 -41004 3100
rect -34825 -3100 -34765 3100
rect -34745 -3100 -34685 3100
rect -28506 -3100 -28446 3100
rect -28426 -3100 -28366 3100
rect -22187 -3100 -22127 3100
rect -22107 -3100 -22047 3100
rect -15868 -3100 -15808 3100
rect -15788 -3100 -15728 3100
rect -9549 -3100 -9489 3100
rect -9469 -3100 -9409 3100
rect -3230 -3100 -3170 3100
rect -3150 -3100 -3090 3100
rect 3089 -3100 3149 3100
rect 3169 -3100 3229 3100
rect 9408 -3100 9468 3100
rect 9488 -3100 9548 3100
rect 15727 -3100 15787 3100
rect 15807 -3100 15867 3100
rect 22046 -3100 22106 3100
rect 22126 -3100 22186 3100
rect 28365 -3100 28425 3100
rect 28445 -3100 28505 3100
rect 34684 -3100 34744 3100
rect 34764 -3100 34824 3100
rect 41003 -3100 41063 3100
rect 41083 -3100 41143 3100
rect -41144 -9400 -41084 -3200
rect -41064 -9400 -41004 -3200
rect -34825 -9400 -34765 -3200
rect -34745 -9400 -34685 -3200
rect -28506 -9400 -28446 -3200
rect -28426 -9400 -28366 -3200
rect -22187 -9400 -22127 -3200
rect -22107 -9400 -22047 -3200
rect -15868 -9400 -15808 -3200
rect -15788 -9400 -15728 -3200
rect -9549 -9400 -9489 -3200
rect -9469 -9400 -9409 -3200
rect -3230 -9400 -3170 -3200
rect -3150 -9400 -3090 -3200
rect 3089 -9400 3149 -3200
rect 3169 -9400 3229 -3200
rect 9408 -9400 9468 -3200
rect 9488 -9400 9548 -3200
rect 15727 -9400 15787 -3200
rect 15807 -9400 15867 -3200
rect 22046 -9400 22106 -3200
rect 22126 -9400 22186 -3200
rect 28365 -9400 28425 -3200
rect 28445 -9400 28505 -3200
rect 34684 -9400 34744 -3200
rect 34764 -9400 34824 -3200
rect 41003 -9400 41063 -3200
rect 41083 -9400 41143 -3200
rect -41144 -15700 -41084 -9500
rect -41064 -15700 -41004 -9500
rect -34825 -15700 -34765 -9500
rect -34745 -15700 -34685 -9500
rect -28506 -15700 -28446 -9500
rect -28426 -15700 -28366 -9500
rect -22187 -15700 -22127 -9500
rect -22107 -15700 -22047 -9500
rect -15868 -15700 -15808 -9500
rect -15788 -15700 -15728 -9500
rect -9549 -15700 -9489 -9500
rect -9469 -15700 -9409 -9500
rect -3230 -15700 -3170 -9500
rect -3150 -15700 -3090 -9500
rect 3089 -15700 3149 -9500
rect 3169 -15700 3229 -9500
rect 9408 -15700 9468 -9500
rect 9488 -15700 9548 -9500
rect 15727 -15700 15787 -9500
rect 15807 -15700 15867 -9500
rect 22046 -15700 22106 -9500
rect 22126 -15700 22186 -9500
rect 28365 -15700 28425 -9500
rect 28445 -15700 28505 -9500
rect 34684 -15700 34744 -9500
rect 34764 -15700 34824 -9500
rect 41003 -15700 41063 -9500
rect 41083 -15700 41143 -9500
rect -41144 -22000 -41084 -15800
rect -41064 -22000 -41004 -15800
rect -34825 -22000 -34765 -15800
rect -34745 -22000 -34685 -15800
rect -28506 -22000 -28446 -15800
rect -28426 -22000 -28366 -15800
rect -22187 -22000 -22127 -15800
rect -22107 -22000 -22047 -15800
rect -15868 -22000 -15808 -15800
rect -15788 -22000 -15728 -15800
rect -9549 -22000 -9489 -15800
rect -9469 -22000 -9409 -15800
rect -3230 -22000 -3170 -15800
rect -3150 -22000 -3090 -15800
rect 3089 -22000 3149 -15800
rect 3169 -22000 3229 -15800
rect 9408 -22000 9468 -15800
rect 9488 -22000 9548 -15800
rect 15727 -22000 15787 -15800
rect 15807 -22000 15867 -15800
rect 22046 -22000 22106 -15800
rect 22126 -22000 22186 -15800
rect 28365 -22000 28425 -15800
rect 28445 -22000 28505 -15800
rect 34684 -22000 34744 -15800
rect 34764 -22000 34824 -15800
rect 41003 -22000 41063 -15800
rect 41083 -22000 41143 -15800
rect -41144 -28300 -41084 -22100
rect -41064 -28300 -41004 -22100
rect -34825 -28300 -34765 -22100
rect -34745 -28300 -34685 -22100
rect -28506 -28300 -28446 -22100
rect -28426 -28300 -28366 -22100
rect -22187 -28300 -22127 -22100
rect -22107 -28300 -22047 -22100
rect -15868 -28300 -15808 -22100
rect -15788 -28300 -15728 -22100
rect -9549 -28300 -9489 -22100
rect -9469 -28300 -9409 -22100
rect -3230 -28300 -3170 -22100
rect -3150 -28300 -3090 -22100
rect 3089 -28300 3149 -22100
rect 3169 -28300 3229 -22100
rect 9408 -28300 9468 -22100
rect 9488 -28300 9548 -22100
rect 15727 -28300 15787 -22100
rect 15807 -28300 15867 -22100
rect 22046 -28300 22106 -22100
rect 22126 -28300 22186 -22100
rect 28365 -28300 28425 -22100
rect 28445 -28300 28505 -22100
rect 34684 -28300 34744 -22100
rect 34764 -28300 34824 -22100
rect 41003 -28300 41063 -22100
rect 41083 -28300 41143 -22100
rect -41144 -34600 -41084 -28400
rect -41064 -34600 -41004 -28400
rect -34825 -34600 -34765 -28400
rect -34745 -34600 -34685 -28400
rect -28506 -34600 -28446 -28400
rect -28426 -34600 -28366 -28400
rect -22187 -34600 -22127 -28400
rect -22107 -34600 -22047 -28400
rect -15868 -34600 -15808 -28400
rect -15788 -34600 -15728 -28400
rect -9549 -34600 -9489 -28400
rect -9469 -34600 -9409 -28400
rect -3230 -34600 -3170 -28400
rect -3150 -34600 -3090 -28400
rect 3089 -34600 3149 -28400
rect 3169 -34600 3229 -28400
rect 9408 -34600 9468 -28400
rect 9488 -34600 9548 -28400
rect 15727 -34600 15787 -28400
rect 15807 -34600 15867 -28400
rect 22046 -34600 22106 -28400
rect 22126 -34600 22186 -28400
rect 28365 -34600 28425 -28400
rect 28445 -34600 28505 -28400
rect 34684 -34600 34744 -28400
rect 34764 -34600 34824 -28400
rect 41003 -34600 41063 -28400
rect 41083 -34600 41143 -28400
rect -41144 -40900 -41084 -34700
rect -41064 -40900 -41004 -34700
rect -34825 -40900 -34765 -34700
rect -34745 -40900 -34685 -34700
rect -28506 -40900 -28446 -34700
rect -28426 -40900 -28366 -34700
rect -22187 -40900 -22127 -34700
rect -22107 -40900 -22047 -34700
rect -15868 -40900 -15808 -34700
rect -15788 -40900 -15728 -34700
rect -9549 -40900 -9489 -34700
rect -9469 -40900 -9409 -34700
rect -3230 -40900 -3170 -34700
rect -3150 -40900 -3090 -34700
rect 3089 -40900 3149 -34700
rect 3169 -40900 3229 -34700
rect 9408 -40900 9468 -34700
rect 9488 -40900 9548 -34700
rect 15727 -40900 15787 -34700
rect 15807 -40900 15867 -34700
rect 22046 -40900 22106 -34700
rect 22126 -40900 22186 -34700
rect 28365 -40900 28425 -34700
rect 28445 -40900 28505 -34700
rect 34684 -40900 34744 -34700
rect 34764 -40900 34824 -34700
rect 41003 -40900 41063 -34700
rect 41083 -40900 41143 -34700
rect -41144 -47200 -41084 -41000
rect -41064 -47200 -41004 -41000
rect -34825 -47200 -34765 -41000
rect -34745 -47200 -34685 -41000
rect -28506 -47200 -28446 -41000
rect -28426 -47200 -28366 -41000
rect -22187 -47200 -22127 -41000
rect -22107 -47200 -22047 -41000
rect -15868 -47200 -15808 -41000
rect -15788 -47200 -15728 -41000
rect -9549 -47200 -9489 -41000
rect -9469 -47200 -9409 -41000
rect -3230 -47200 -3170 -41000
rect -3150 -47200 -3090 -41000
rect 3089 -47200 3149 -41000
rect 3169 -47200 3229 -41000
rect 9408 -47200 9468 -41000
rect 9488 -47200 9548 -41000
rect 15727 -47200 15787 -41000
rect 15807 -47200 15867 -41000
rect 22046 -47200 22106 -41000
rect 22126 -47200 22186 -41000
rect 28365 -47200 28425 -41000
rect 28445 -47200 28505 -41000
rect 34684 -47200 34744 -41000
rect 34764 -47200 34824 -41000
rect 41003 -47200 41063 -41000
rect 41083 -47200 41143 -41000
<< metal3 >>
rect -47383 47172 -41084 47200
rect -47383 41028 -41168 47172
rect -41104 41028 -41084 47172
rect -47383 41000 -41084 41028
rect -41064 47172 -34765 47200
rect -41064 41028 -34849 47172
rect -34785 41028 -34765 47172
rect -41064 41000 -34765 41028
rect -34745 47172 -28446 47200
rect -34745 41028 -28530 47172
rect -28466 41028 -28446 47172
rect -34745 41000 -28446 41028
rect -28426 47172 -22127 47200
rect -28426 41028 -22211 47172
rect -22147 41028 -22127 47172
rect -28426 41000 -22127 41028
rect -22107 47172 -15808 47200
rect -22107 41028 -15892 47172
rect -15828 41028 -15808 47172
rect -22107 41000 -15808 41028
rect -15788 47172 -9489 47200
rect -15788 41028 -9573 47172
rect -9509 41028 -9489 47172
rect -15788 41000 -9489 41028
rect -9469 47172 -3170 47200
rect -9469 41028 -3254 47172
rect -3190 41028 -3170 47172
rect -9469 41000 -3170 41028
rect -3150 47172 3149 47200
rect -3150 41028 3065 47172
rect 3129 41028 3149 47172
rect -3150 41000 3149 41028
rect 3169 47172 9468 47200
rect 3169 41028 9384 47172
rect 9448 41028 9468 47172
rect 3169 41000 9468 41028
rect 9488 47172 15787 47200
rect 9488 41028 15703 47172
rect 15767 41028 15787 47172
rect 9488 41000 15787 41028
rect 15807 47172 22106 47200
rect 15807 41028 22022 47172
rect 22086 41028 22106 47172
rect 15807 41000 22106 41028
rect 22126 47172 28425 47200
rect 22126 41028 28341 47172
rect 28405 41028 28425 47172
rect 22126 41000 28425 41028
rect 28445 47172 34744 47200
rect 28445 41028 34660 47172
rect 34724 41028 34744 47172
rect 28445 41000 34744 41028
rect 34764 47172 41063 47200
rect 34764 41028 40979 47172
rect 41043 41028 41063 47172
rect 34764 41000 41063 41028
rect 41083 47172 47382 47200
rect 41083 41028 47298 47172
rect 47362 41028 47382 47172
rect 41083 41000 47382 41028
rect -47383 40872 -41084 40900
rect -47383 34728 -41168 40872
rect -41104 34728 -41084 40872
rect -47383 34700 -41084 34728
rect -41064 40872 -34765 40900
rect -41064 34728 -34849 40872
rect -34785 34728 -34765 40872
rect -41064 34700 -34765 34728
rect -34745 40872 -28446 40900
rect -34745 34728 -28530 40872
rect -28466 34728 -28446 40872
rect -34745 34700 -28446 34728
rect -28426 40872 -22127 40900
rect -28426 34728 -22211 40872
rect -22147 34728 -22127 40872
rect -28426 34700 -22127 34728
rect -22107 40872 -15808 40900
rect -22107 34728 -15892 40872
rect -15828 34728 -15808 40872
rect -22107 34700 -15808 34728
rect -15788 40872 -9489 40900
rect -15788 34728 -9573 40872
rect -9509 34728 -9489 40872
rect -15788 34700 -9489 34728
rect -9469 40872 -3170 40900
rect -9469 34728 -3254 40872
rect -3190 34728 -3170 40872
rect -9469 34700 -3170 34728
rect -3150 40872 3149 40900
rect -3150 34728 3065 40872
rect 3129 34728 3149 40872
rect -3150 34700 3149 34728
rect 3169 40872 9468 40900
rect 3169 34728 9384 40872
rect 9448 34728 9468 40872
rect 3169 34700 9468 34728
rect 9488 40872 15787 40900
rect 9488 34728 15703 40872
rect 15767 34728 15787 40872
rect 9488 34700 15787 34728
rect 15807 40872 22106 40900
rect 15807 34728 22022 40872
rect 22086 34728 22106 40872
rect 15807 34700 22106 34728
rect 22126 40872 28425 40900
rect 22126 34728 28341 40872
rect 28405 34728 28425 40872
rect 22126 34700 28425 34728
rect 28445 40872 34744 40900
rect 28445 34728 34660 40872
rect 34724 34728 34744 40872
rect 28445 34700 34744 34728
rect 34764 40872 41063 40900
rect 34764 34728 40979 40872
rect 41043 34728 41063 40872
rect 34764 34700 41063 34728
rect 41083 40872 47382 40900
rect 41083 34728 47298 40872
rect 47362 34728 47382 40872
rect 41083 34700 47382 34728
rect -47383 34572 -41084 34600
rect -47383 28428 -41168 34572
rect -41104 28428 -41084 34572
rect -47383 28400 -41084 28428
rect -41064 34572 -34765 34600
rect -41064 28428 -34849 34572
rect -34785 28428 -34765 34572
rect -41064 28400 -34765 28428
rect -34745 34572 -28446 34600
rect -34745 28428 -28530 34572
rect -28466 28428 -28446 34572
rect -34745 28400 -28446 28428
rect -28426 34572 -22127 34600
rect -28426 28428 -22211 34572
rect -22147 28428 -22127 34572
rect -28426 28400 -22127 28428
rect -22107 34572 -15808 34600
rect -22107 28428 -15892 34572
rect -15828 28428 -15808 34572
rect -22107 28400 -15808 28428
rect -15788 34572 -9489 34600
rect -15788 28428 -9573 34572
rect -9509 28428 -9489 34572
rect -15788 28400 -9489 28428
rect -9469 34572 -3170 34600
rect -9469 28428 -3254 34572
rect -3190 28428 -3170 34572
rect -9469 28400 -3170 28428
rect -3150 34572 3149 34600
rect -3150 28428 3065 34572
rect 3129 28428 3149 34572
rect -3150 28400 3149 28428
rect 3169 34572 9468 34600
rect 3169 28428 9384 34572
rect 9448 28428 9468 34572
rect 3169 28400 9468 28428
rect 9488 34572 15787 34600
rect 9488 28428 15703 34572
rect 15767 28428 15787 34572
rect 9488 28400 15787 28428
rect 15807 34572 22106 34600
rect 15807 28428 22022 34572
rect 22086 28428 22106 34572
rect 15807 28400 22106 28428
rect 22126 34572 28425 34600
rect 22126 28428 28341 34572
rect 28405 28428 28425 34572
rect 22126 28400 28425 28428
rect 28445 34572 34744 34600
rect 28445 28428 34660 34572
rect 34724 28428 34744 34572
rect 28445 28400 34744 28428
rect 34764 34572 41063 34600
rect 34764 28428 40979 34572
rect 41043 28428 41063 34572
rect 34764 28400 41063 28428
rect 41083 34572 47382 34600
rect 41083 28428 47298 34572
rect 47362 28428 47382 34572
rect 41083 28400 47382 28428
rect -47383 28272 -41084 28300
rect -47383 22128 -41168 28272
rect -41104 22128 -41084 28272
rect -47383 22100 -41084 22128
rect -41064 28272 -34765 28300
rect -41064 22128 -34849 28272
rect -34785 22128 -34765 28272
rect -41064 22100 -34765 22128
rect -34745 28272 -28446 28300
rect -34745 22128 -28530 28272
rect -28466 22128 -28446 28272
rect -34745 22100 -28446 22128
rect -28426 28272 -22127 28300
rect -28426 22128 -22211 28272
rect -22147 22128 -22127 28272
rect -28426 22100 -22127 22128
rect -22107 28272 -15808 28300
rect -22107 22128 -15892 28272
rect -15828 22128 -15808 28272
rect -22107 22100 -15808 22128
rect -15788 28272 -9489 28300
rect -15788 22128 -9573 28272
rect -9509 22128 -9489 28272
rect -15788 22100 -9489 22128
rect -9469 28272 -3170 28300
rect -9469 22128 -3254 28272
rect -3190 22128 -3170 28272
rect -9469 22100 -3170 22128
rect -3150 28272 3149 28300
rect -3150 22128 3065 28272
rect 3129 22128 3149 28272
rect -3150 22100 3149 22128
rect 3169 28272 9468 28300
rect 3169 22128 9384 28272
rect 9448 22128 9468 28272
rect 3169 22100 9468 22128
rect 9488 28272 15787 28300
rect 9488 22128 15703 28272
rect 15767 22128 15787 28272
rect 9488 22100 15787 22128
rect 15807 28272 22106 28300
rect 15807 22128 22022 28272
rect 22086 22128 22106 28272
rect 15807 22100 22106 22128
rect 22126 28272 28425 28300
rect 22126 22128 28341 28272
rect 28405 22128 28425 28272
rect 22126 22100 28425 22128
rect 28445 28272 34744 28300
rect 28445 22128 34660 28272
rect 34724 22128 34744 28272
rect 28445 22100 34744 22128
rect 34764 28272 41063 28300
rect 34764 22128 40979 28272
rect 41043 22128 41063 28272
rect 34764 22100 41063 22128
rect 41083 28272 47382 28300
rect 41083 22128 47298 28272
rect 47362 22128 47382 28272
rect 41083 22100 47382 22128
rect -47383 21972 -41084 22000
rect -47383 15828 -41168 21972
rect -41104 15828 -41084 21972
rect -47383 15800 -41084 15828
rect -41064 21972 -34765 22000
rect -41064 15828 -34849 21972
rect -34785 15828 -34765 21972
rect -41064 15800 -34765 15828
rect -34745 21972 -28446 22000
rect -34745 15828 -28530 21972
rect -28466 15828 -28446 21972
rect -34745 15800 -28446 15828
rect -28426 21972 -22127 22000
rect -28426 15828 -22211 21972
rect -22147 15828 -22127 21972
rect -28426 15800 -22127 15828
rect -22107 21972 -15808 22000
rect -22107 15828 -15892 21972
rect -15828 15828 -15808 21972
rect -22107 15800 -15808 15828
rect -15788 21972 -9489 22000
rect -15788 15828 -9573 21972
rect -9509 15828 -9489 21972
rect -15788 15800 -9489 15828
rect -9469 21972 -3170 22000
rect -9469 15828 -3254 21972
rect -3190 15828 -3170 21972
rect -9469 15800 -3170 15828
rect -3150 21972 3149 22000
rect -3150 15828 3065 21972
rect 3129 15828 3149 21972
rect -3150 15800 3149 15828
rect 3169 21972 9468 22000
rect 3169 15828 9384 21972
rect 9448 15828 9468 21972
rect 3169 15800 9468 15828
rect 9488 21972 15787 22000
rect 9488 15828 15703 21972
rect 15767 15828 15787 21972
rect 9488 15800 15787 15828
rect 15807 21972 22106 22000
rect 15807 15828 22022 21972
rect 22086 15828 22106 21972
rect 15807 15800 22106 15828
rect 22126 21972 28425 22000
rect 22126 15828 28341 21972
rect 28405 15828 28425 21972
rect 22126 15800 28425 15828
rect 28445 21972 34744 22000
rect 28445 15828 34660 21972
rect 34724 15828 34744 21972
rect 28445 15800 34744 15828
rect 34764 21972 41063 22000
rect 34764 15828 40979 21972
rect 41043 15828 41063 21972
rect 34764 15800 41063 15828
rect 41083 21972 47382 22000
rect 41083 15828 47298 21972
rect 47362 15828 47382 21972
rect 41083 15800 47382 15828
rect -47383 15672 -41084 15700
rect -47383 9528 -41168 15672
rect -41104 9528 -41084 15672
rect -47383 9500 -41084 9528
rect -41064 15672 -34765 15700
rect -41064 9528 -34849 15672
rect -34785 9528 -34765 15672
rect -41064 9500 -34765 9528
rect -34745 15672 -28446 15700
rect -34745 9528 -28530 15672
rect -28466 9528 -28446 15672
rect -34745 9500 -28446 9528
rect -28426 15672 -22127 15700
rect -28426 9528 -22211 15672
rect -22147 9528 -22127 15672
rect -28426 9500 -22127 9528
rect -22107 15672 -15808 15700
rect -22107 9528 -15892 15672
rect -15828 9528 -15808 15672
rect -22107 9500 -15808 9528
rect -15788 15672 -9489 15700
rect -15788 9528 -9573 15672
rect -9509 9528 -9489 15672
rect -15788 9500 -9489 9528
rect -9469 15672 -3170 15700
rect -9469 9528 -3254 15672
rect -3190 9528 -3170 15672
rect -9469 9500 -3170 9528
rect -3150 15672 3149 15700
rect -3150 9528 3065 15672
rect 3129 9528 3149 15672
rect -3150 9500 3149 9528
rect 3169 15672 9468 15700
rect 3169 9528 9384 15672
rect 9448 9528 9468 15672
rect 3169 9500 9468 9528
rect 9488 15672 15787 15700
rect 9488 9528 15703 15672
rect 15767 9528 15787 15672
rect 9488 9500 15787 9528
rect 15807 15672 22106 15700
rect 15807 9528 22022 15672
rect 22086 9528 22106 15672
rect 15807 9500 22106 9528
rect 22126 15672 28425 15700
rect 22126 9528 28341 15672
rect 28405 9528 28425 15672
rect 22126 9500 28425 9528
rect 28445 15672 34744 15700
rect 28445 9528 34660 15672
rect 34724 9528 34744 15672
rect 28445 9500 34744 9528
rect 34764 15672 41063 15700
rect 34764 9528 40979 15672
rect 41043 9528 41063 15672
rect 34764 9500 41063 9528
rect 41083 15672 47382 15700
rect 41083 9528 47298 15672
rect 47362 9528 47382 15672
rect 41083 9500 47382 9528
rect -47383 9372 -41084 9400
rect -47383 3228 -41168 9372
rect -41104 3228 -41084 9372
rect -47383 3200 -41084 3228
rect -41064 9372 -34765 9400
rect -41064 3228 -34849 9372
rect -34785 3228 -34765 9372
rect -41064 3200 -34765 3228
rect -34745 9372 -28446 9400
rect -34745 3228 -28530 9372
rect -28466 3228 -28446 9372
rect -34745 3200 -28446 3228
rect -28426 9372 -22127 9400
rect -28426 3228 -22211 9372
rect -22147 3228 -22127 9372
rect -28426 3200 -22127 3228
rect -22107 9372 -15808 9400
rect -22107 3228 -15892 9372
rect -15828 3228 -15808 9372
rect -22107 3200 -15808 3228
rect -15788 9372 -9489 9400
rect -15788 3228 -9573 9372
rect -9509 3228 -9489 9372
rect -15788 3200 -9489 3228
rect -9469 9372 -3170 9400
rect -9469 3228 -3254 9372
rect -3190 3228 -3170 9372
rect -9469 3200 -3170 3228
rect -3150 9372 3149 9400
rect -3150 3228 3065 9372
rect 3129 3228 3149 9372
rect -3150 3200 3149 3228
rect 3169 9372 9468 9400
rect 3169 3228 9384 9372
rect 9448 3228 9468 9372
rect 3169 3200 9468 3228
rect 9488 9372 15787 9400
rect 9488 3228 15703 9372
rect 15767 3228 15787 9372
rect 9488 3200 15787 3228
rect 15807 9372 22106 9400
rect 15807 3228 22022 9372
rect 22086 3228 22106 9372
rect 15807 3200 22106 3228
rect 22126 9372 28425 9400
rect 22126 3228 28341 9372
rect 28405 3228 28425 9372
rect 22126 3200 28425 3228
rect 28445 9372 34744 9400
rect 28445 3228 34660 9372
rect 34724 3228 34744 9372
rect 28445 3200 34744 3228
rect 34764 9372 41063 9400
rect 34764 3228 40979 9372
rect 41043 3228 41063 9372
rect 34764 3200 41063 3228
rect 41083 9372 47382 9400
rect 41083 3228 47298 9372
rect 47362 3228 47382 9372
rect 41083 3200 47382 3228
rect -47383 3072 -41084 3100
rect -47383 -3072 -41168 3072
rect -41104 -3072 -41084 3072
rect -47383 -3100 -41084 -3072
rect -41064 3072 -34765 3100
rect -41064 -3072 -34849 3072
rect -34785 -3072 -34765 3072
rect -41064 -3100 -34765 -3072
rect -34745 3072 -28446 3100
rect -34745 -3072 -28530 3072
rect -28466 -3072 -28446 3072
rect -34745 -3100 -28446 -3072
rect -28426 3072 -22127 3100
rect -28426 -3072 -22211 3072
rect -22147 -3072 -22127 3072
rect -28426 -3100 -22127 -3072
rect -22107 3072 -15808 3100
rect -22107 -3072 -15892 3072
rect -15828 -3072 -15808 3072
rect -22107 -3100 -15808 -3072
rect -15788 3072 -9489 3100
rect -15788 -3072 -9573 3072
rect -9509 -3072 -9489 3072
rect -15788 -3100 -9489 -3072
rect -9469 3072 -3170 3100
rect -9469 -3072 -3254 3072
rect -3190 -3072 -3170 3072
rect -9469 -3100 -3170 -3072
rect -3150 3072 3149 3100
rect -3150 -3072 3065 3072
rect 3129 -3072 3149 3072
rect -3150 -3100 3149 -3072
rect 3169 3072 9468 3100
rect 3169 -3072 9384 3072
rect 9448 -3072 9468 3072
rect 3169 -3100 9468 -3072
rect 9488 3072 15787 3100
rect 9488 -3072 15703 3072
rect 15767 -3072 15787 3072
rect 9488 -3100 15787 -3072
rect 15807 3072 22106 3100
rect 15807 -3072 22022 3072
rect 22086 -3072 22106 3072
rect 15807 -3100 22106 -3072
rect 22126 3072 28425 3100
rect 22126 -3072 28341 3072
rect 28405 -3072 28425 3072
rect 22126 -3100 28425 -3072
rect 28445 3072 34744 3100
rect 28445 -3072 34660 3072
rect 34724 -3072 34744 3072
rect 28445 -3100 34744 -3072
rect 34764 3072 41063 3100
rect 34764 -3072 40979 3072
rect 41043 -3072 41063 3072
rect 34764 -3100 41063 -3072
rect 41083 3072 47382 3100
rect 41083 -3072 47298 3072
rect 47362 -3072 47382 3072
rect 41083 -3100 47382 -3072
rect -47383 -3228 -41084 -3200
rect -47383 -9372 -41168 -3228
rect -41104 -9372 -41084 -3228
rect -47383 -9400 -41084 -9372
rect -41064 -3228 -34765 -3200
rect -41064 -9372 -34849 -3228
rect -34785 -9372 -34765 -3228
rect -41064 -9400 -34765 -9372
rect -34745 -3228 -28446 -3200
rect -34745 -9372 -28530 -3228
rect -28466 -9372 -28446 -3228
rect -34745 -9400 -28446 -9372
rect -28426 -3228 -22127 -3200
rect -28426 -9372 -22211 -3228
rect -22147 -9372 -22127 -3228
rect -28426 -9400 -22127 -9372
rect -22107 -3228 -15808 -3200
rect -22107 -9372 -15892 -3228
rect -15828 -9372 -15808 -3228
rect -22107 -9400 -15808 -9372
rect -15788 -3228 -9489 -3200
rect -15788 -9372 -9573 -3228
rect -9509 -9372 -9489 -3228
rect -15788 -9400 -9489 -9372
rect -9469 -3228 -3170 -3200
rect -9469 -9372 -3254 -3228
rect -3190 -9372 -3170 -3228
rect -9469 -9400 -3170 -9372
rect -3150 -3228 3149 -3200
rect -3150 -9372 3065 -3228
rect 3129 -9372 3149 -3228
rect -3150 -9400 3149 -9372
rect 3169 -3228 9468 -3200
rect 3169 -9372 9384 -3228
rect 9448 -9372 9468 -3228
rect 3169 -9400 9468 -9372
rect 9488 -3228 15787 -3200
rect 9488 -9372 15703 -3228
rect 15767 -9372 15787 -3228
rect 9488 -9400 15787 -9372
rect 15807 -3228 22106 -3200
rect 15807 -9372 22022 -3228
rect 22086 -9372 22106 -3228
rect 15807 -9400 22106 -9372
rect 22126 -3228 28425 -3200
rect 22126 -9372 28341 -3228
rect 28405 -9372 28425 -3228
rect 22126 -9400 28425 -9372
rect 28445 -3228 34744 -3200
rect 28445 -9372 34660 -3228
rect 34724 -9372 34744 -3228
rect 28445 -9400 34744 -9372
rect 34764 -3228 41063 -3200
rect 34764 -9372 40979 -3228
rect 41043 -9372 41063 -3228
rect 34764 -9400 41063 -9372
rect 41083 -3228 47382 -3200
rect 41083 -9372 47298 -3228
rect 47362 -9372 47382 -3228
rect 41083 -9400 47382 -9372
rect -47383 -9528 -41084 -9500
rect -47383 -15672 -41168 -9528
rect -41104 -15672 -41084 -9528
rect -47383 -15700 -41084 -15672
rect -41064 -9528 -34765 -9500
rect -41064 -15672 -34849 -9528
rect -34785 -15672 -34765 -9528
rect -41064 -15700 -34765 -15672
rect -34745 -9528 -28446 -9500
rect -34745 -15672 -28530 -9528
rect -28466 -15672 -28446 -9528
rect -34745 -15700 -28446 -15672
rect -28426 -9528 -22127 -9500
rect -28426 -15672 -22211 -9528
rect -22147 -15672 -22127 -9528
rect -28426 -15700 -22127 -15672
rect -22107 -9528 -15808 -9500
rect -22107 -15672 -15892 -9528
rect -15828 -15672 -15808 -9528
rect -22107 -15700 -15808 -15672
rect -15788 -9528 -9489 -9500
rect -15788 -15672 -9573 -9528
rect -9509 -15672 -9489 -9528
rect -15788 -15700 -9489 -15672
rect -9469 -9528 -3170 -9500
rect -9469 -15672 -3254 -9528
rect -3190 -15672 -3170 -9528
rect -9469 -15700 -3170 -15672
rect -3150 -9528 3149 -9500
rect -3150 -15672 3065 -9528
rect 3129 -15672 3149 -9528
rect -3150 -15700 3149 -15672
rect 3169 -9528 9468 -9500
rect 3169 -15672 9384 -9528
rect 9448 -15672 9468 -9528
rect 3169 -15700 9468 -15672
rect 9488 -9528 15787 -9500
rect 9488 -15672 15703 -9528
rect 15767 -15672 15787 -9528
rect 9488 -15700 15787 -15672
rect 15807 -9528 22106 -9500
rect 15807 -15672 22022 -9528
rect 22086 -15672 22106 -9528
rect 15807 -15700 22106 -15672
rect 22126 -9528 28425 -9500
rect 22126 -15672 28341 -9528
rect 28405 -15672 28425 -9528
rect 22126 -15700 28425 -15672
rect 28445 -9528 34744 -9500
rect 28445 -15672 34660 -9528
rect 34724 -15672 34744 -9528
rect 28445 -15700 34744 -15672
rect 34764 -9528 41063 -9500
rect 34764 -15672 40979 -9528
rect 41043 -15672 41063 -9528
rect 34764 -15700 41063 -15672
rect 41083 -9528 47382 -9500
rect 41083 -15672 47298 -9528
rect 47362 -15672 47382 -9528
rect 41083 -15700 47382 -15672
rect -47383 -15828 -41084 -15800
rect -47383 -21972 -41168 -15828
rect -41104 -21972 -41084 -15828
rect -47383 -22000 -41084 -21972
rect -41064 -15828 -34765 -15800
rect -41064 -21972 -34849 -15828
rect -34785 -21972 -34765 -15828
rect -41064 -22000 -34765 -21972
rect -34745 -15828 -28446 -15800
rect -34745 -21972 -28530 -15828
rect -28466 -21972 -28446 -15828
rect -34745 -22000 -28446 -21972
rect -28426 -15828 -22127 -15800
rect -28426 -21972 -22211 -15828
rect -22147 -21972 -22127 -15828
rect -28426 -22000 -22127 -21972
rect -22107 -15828 -15808 -15800
rect -22107 -21972 -15892 -15828
rect -15828 -21972 -15808 -15828
rect -22107 -22000 -15808 -21972
rect -15788 -15828 -9489 -15800
rect -15788 -21972 -9573 -15828
rect -9509 -21972 -9489 -15828
rect -15788 -22000 -9489 -21972
rect -9469 -15828 -3170 -15800
rect -9469 -21972 -3254 -15828
rect -3190 -21972 -3170 -15828
rect -9469 -22000 -3170 -21972
rect -3150 -15828 3149 -15800
rect -3150 -21972 3065 -15828
rect 3129 -21972 3149 -15828
rect -3150 -22000 3149 -21972
rect 3169 -15828 9468 -15800
rect 3169 -21972 9384 -15828
rect 9448 -21972 9468 -15828
rect 3169 -22000 9468 -21972
rect 9488 -15828 15787 -15800
rect 9488 -21972 15703 -15828
rect 15767 -21972 15787 -15828
rect 9488 -22000 15787 -21972
rect 15807 -15828 22106 -15800
rect 15807 -21972 22022 -15828
rect 22086 -21972 22106 -15828
rect 15807 -22000 22106 -21972
rect 22126 -15828 28425 -15800
rect 22126 -21972 28341 -15828
rect 28405 -21972 28425 -15828
rect 22126 -22000 28425 -21972
rect 28445 -15828 34744 -15800
rect 28445 -21972 34660 -15828
rect 34724 -21972 34744 -15828
rect 28445 -22000 34744 -21972
rect 34764 -15828 41063 -15800
rect 34764 -21972 40979 -15828
rect 41043 -21972 41063 -15828
rect 34764 -22000 41063 -21972
rect 41083 -15828 47382 -15800
rect 41083 -21972 47298 -15828
rect 47362 -21972 47382 -15828
rect 41083 -22000 47382 -21972
rect -47383 -22128 -41084 -22100
rect -47383 -28272 -41168 -22128
rect -41104 -28272 -41084 -22128
rect -47383 -28300 -41084 -28272
rect -41064 -22128 -34765 -22100
rect -41064 -28272 -34849 -22128
rect -34785 -28272 -34765 -22128
rect -41064 -28300 -34765 -28272
rect -34745 -22128 -28446 -22100
rect -34745 -28272 -28530 -22128
rect -28466 -28272 -28446 -22128
rect -34745 -28300 -28446 -28272
rect -28426 -22128 -22127 -22100
rect -28426 -28272 -22211 -22128
rect -22147 -28272 -22127 -22128
rect -28426 -28300 -22127 -28272
rect -22107 -22128 -15808 -22100
rect -22107 -28272 -15892 -22128
rect -15828 -28272 -15808 -22128
rect -22107 -28300 -15808 -28272
rect -15788 -22128 -9489 -22100
rect -15788 -28272 -9573 -22128
rect -9509 -28272 -9489 -22128
rect -15788 -28300 -9489 -28272
rect -9469 -22128 -3170 -22100
rect -9469 -28272 -3254 -22128
rect -3190 -28272 -3170 -22128
rect -9469 -28300 -3170 -28272
rect -3150 -22128 3149 -22100
rect -3150 -28272 3065 -22128
rect 3129 -28272 3149 -22128
rect -3150 -28300 3149 -28272
rect 3169 -22128 9468 -22100
rect 3169 -28272 9384 -22128
rect 9448 -28272 9468 -22128
rect 3169 -28300 9468 -28272
rect 9488 -22128 15787 -22100
rect 9488 -28272 15703 -22128
rect 15767 -28272 15787 -22128
rect 9488 -28300 15787 -28272
rect 15807 -22128 22106 -22100
rect 15807 -28272 22022 -22128
rect 22086 -28272 22106 -22128
rect 15807 -28300 22106 -28272
rect 22126 -22128 28425 -22100
rect 22126 -28272 28341 -22128
rect 28405 -28272 28425 -22128
rect 22126 -28300 28425 -28272
rect 28445 -22128 34744 -22100
rect 28445 -28272 34660 -22128
rect 34724 -28272 34744 -22128
rect 28445 -28300 34744 -28272
rect 34764 -22128 41063 -22100
rect 34764 -28272 40979 -22128
rect 41043 -28272 41063 -22128
rect 34764 -28300 41063 -28272
rect 41083 -22128 47382 -22100
rect 41083 -28272 47298 -22128
rect 47362 -28272 47382 -22128
rect 41083 -28300 47382 -28272
rect -47383 -28428 -41084 -28400
rect -47383 -34572 -41168 -28428
rect -41104 -34572 -41084 -28428
rect -47383 -34600 -41084 -34572
rect -41064 -28428 -34765 -28400
rect -41064 -34572 -34849 -28428
rect -34785 -34572 -34765 -28428
rect -41064 -34600 -34765 -34572
rect -34745 -28428 -28446 -28400
rect -34745 -34572 -28530 -28428
rect -28466 -34572 -28446 -28428
rect -34745 -34600 -28446 -34572
rect -28426 -28428 -22127 -28400
rect -28426 -34572 -22211 -28428
rect -22147 -34572 -22127 -28428
rect -28426 -34600 -22127 -34572
rect -22107 -28428 -15808 -28400
rect -22107 -34572 -15892 -28428
rect -15828 -34572 -15808 -28428
rect -22107 -34600 -15808 -34572
rect -15788 -28428 -9489 -28400
rect -15788 -34572 -9573 -28428
rect -9509 -34572 -9489 -28428
rect -15788 -34600 -9489 -34572
rect -9469 -28428 -3170 -28400
rect -9469 -34572 -3254 -28428
rect -3190 -34572 -3170 -28428
rect -9469 -34600 -3170 -34572
rect -3150 -28428 3149 -28400
rect -3150 -34572 3065 -28428
rect 3129 -34572 3149 -28428
rect -3150 -34600 3149 -34572
rect 3169 -28428 9468 -28400
rect 3169 -34572 9384 -28428
rect 9448 -34572 9468 -28428
rect 3169 -34600 9468 -34572
rect 9488 -28428 15787 -28400
rect 9488 -34572 15703 -28428
rect 15767 -34572 15787 -28428
rect 9488 -34600 15787 -34572
rect 15807 -28428 22106 -28400
rect 15807 -34572 22022 -28428
rect 22086 -34572 22106 -28428
rect 15807 -34600 22106 -34572
rect 22126 -28428 28425 -28400
rect 22126 -34572 28341 -28428
rect 28405 -34572 28425 -28428
rect 22126 -34600 28425 -34572
rect 28445 -28428 34744 -28400
rect 28445 -34572 34660 -28428
rect 34724 -34572 34744 -28428
rect 28445 -34600 34744 -34572
rect 34764 -28428 41063 -28400
rect 34764 -34572 40979 -28428
rect 41043 -34572 41063 -28428
rect 34764 -34600 41063 -34572
rect 41083 -28428 47382 -28400
rect 41083 -34572 47298 -28428
rect 47362 -34572 47382 -28428
rect 41083 -34600 47382 -34572
rect -47383 -34728 -41084 -34700
rect -47383 -40872 -41168 -34728
rect -41104 -40872 -41084 -34728
rect -47383 -40900 -41084 -40872
rect -41064 -34728 -34765 -34700
rect -41064 -40872 -34849 -34728
rect -34785 -40872 -34765 -34728
rect -41064 -40900 -34765 -40872
rect -34745 -34728 -28446 -34700
rect -34745 -40872 -28530 -34728
rect -28466 -40872 -28446 -34728
rect -34745 -40900 -28446 -40872
rect -28426 -34728 -22127 -34700
rect -28426 -40872 -22211 -34728
rect -22147 -40872 -22127 -34728
rect -28426 -40900 -22127 -40872
rect -22107 -34728 -15808 -34700
rect -22107 -40872 -15892 -34728
rect -15828 -40872 -15808 -34728
rect -22107 -40900 -15808 -40872
rect -15788 -34728 -9489 -34700
rect -15788 -40872 -9573 -34728
rect -9509 -40872 -9489 -34728
rect -15788 -40900 -9489 -40872
rect -9469 -34728 -3170 -34700
rect -9469 -40872 -3254 -34728
rect -3190 -40872 -3170 -34728
rect -9469 -40900 -3170 -40872
rect -3150 -34728 3149 -34700
rect -3150 -40872 3065 -34728
rect 3129 -40872 3149 -34728
rect -3150 -40900 3149 -40872
rect 3169 -34728 9468 -34700
rect 3169 -40872 9384 -34728
rect 9448 -40872 9468 -34728
rect 3169 -40900 9468 -40872
rect 9488 -34728 15787 -34700
rect 9488 -40872 15703 -34728
rect 15767 -40872 15787 -34728
rect 9488 -40900 15787 -40872
rect 15807 -34728 22106 -34700
rect 15807 -40872 22022 -34728
rect 22086 -40872 22106 -34728
rect 15807 -40900 22106 -40872
rect 22126 -34728 28425 -34700
rect 22126 -40872 28341 -34728
rect 28405 -40872 28425 -34728
rect 22126 -40900 28425 -40872
rect 28445 -34728 34744 -34700
rect 28445 -40872 34660 -34728
rect 34724 -40872 34744 -34728
rect 28445 -40900 34744 -40872
rect 34764 -34728 41063 -34700
rect 34764 -40872 40979 -34728
rect 41043 -40872 41063 -34728
rect 34764 -40900 41063 -40872
rect 41083 -34728 47382 -34700
rect 41083 -40872 47298 -34728
rect 47362 -40872 47382 -34728
rect 41083 -40900 47382 -40872
rect -47383 -41028 -41084 -41000
rect -47383 -47172 -41168 -41028
rect -41104 -47172 -41084 -41028
rect -47383 -47200 -41084 -47172
rect -41064 -41028 -34765 -41000
rect -41064 -47172 -34849 -41028
rect -34785 -47172 -34765 -41028
rect -41064 -47200 -34765 -47172
rect -34745 -41028 -28446 -41000
rect -34745 -47172 -28530 -41028
rect -28466 -47172 -28446 -41028
rect -34745 -47200 -28446 -47172
rect -28426 -41028 -22127 -41000
rect -28426 -47172 -22211 -41028
rect -22147 -47172 -22127 -41028
rect -28426 -47200 -22127 -47172
rect -22107 -41028 -15808 -41000
rect -22107 -47172 -15892 -41028
rect -15828 -47172 -15808 -41028
rect -22107 -47200 -15808 -47172
rect -15788 -41028 -9489 -41000
rect -15788 -47172 -9573 -41028
rect -9509 -47172 -9489 -41028
rect -15788 -47200 -9489 -47172
rect -9469 -41028 -3170 -41000
rect -9469 -47172 -3254 -41028
rect -3190 -47172 -3170 -41028
rect -9469 -47200 -3170 -47172
rect -3150 -41028 3149 -41000
rect -3150 -47172 3065 -41028
rect 3129 -47172 3149 -41028
rect -3150 -47200 3149 -47172
rect 3169 -41028 9468 -41000
rect 3169 -47172 9384 -41028
rect 9448 -47172 9468 -41028
rect 3169 -47200 9468 -47172
rect 9488 -41028 15787 -41000
rect 9488 -47172 15703 -41028
rect 15767 -47172 15787 -41028
rect 9488 -47200 15787 -47172
rect 15807 -41028 22106 -41000
rect 15807 -47172 22022 -41028
rect 22086 -47172 22106 -41028
rect 15807 -47200 22106 -47172
rect 22126 -41028 28425 -41000
rect 22126 -47172 28341 -41028
rect 28405 -47172 28425 -41028
rect 22126 -47200 28425 -47172
rect 28445 -41028 34744 -41000
rect 28445 -47172 34660 -41028
rect 34724 -47172 34744 -41028
rect 28445 -47200 34744 -47172
rect 34764 -41028 41063 -41000
rect 34764 -47172 40979 -41028
rect 41043 -47172 41063 -41028
rect 34764 -47200 41063 -47172
rect 41083 -41028 47382 -41000
rect 41083 -47172 47298 -41028
rect 47362 -47172 47382 -41028
rect 41083 -47200 47382 -47172
<< via3 >>
rect -41168 41028 -41104 47172
rect -34849 41028 -34785 47172
rect -28530 41028 -28466 47172
rect -22211 41028 -22147 47172
rect -15892 41028 -15828 47172
rect -9573 41028 -9509 47172
rect -3254 41028 -3190 47172
rect 3065 41028 3129 47172
rect 9384 41028 9448 47172
rect 15703 41028 15767 47172
rect 22022 41028 22086 47172
rect 28341 41028 28405 47172
rect 34660 41028 34724 47172
rect 40979 41028 41043 47172
rect 47298 41028 47362 47172
rect -41168 34728 -41104 40872
rect -34849 34728 -34785 40872
rect -28530 34728 -28466 40872
rect -22211 34728 -22147 40872
rect -15892 34728 -15828 40872
rect -9573 34728 -9509 40872
rect -3254 34728 -3190 40872
rect 3065 34728 3129 40872
rect 9384 34728 9448 40872
rect 15703 34728 15767 40872
rect 22022 34728 22086 40872
rect 28341 34728 28405 40872
rect 34660 34728 34724 40872
rect 40979 34728 41043 40872
rect 47298 34728 47362 40872
rect -41168 28428 -41104 34572
rect -34849 28428 -34785 34572
rect -28530 28428 -28466 34572
rect -22211 28428 -22147 34572
rect -15892 28428 -15828 34572
rect -9573 28428 -9509 34572
rect -3254 28428 -3190 34572
rect 3065 28428 3129 34572
rect 9384 28428 9448 34572
rect 15703 28428 15767 34572
rect 22022 28428 22086 34572
rect 28341 28428 28405 34572
rect 34660 28428 34724 34572
rect 40979 28428 41043 34572
rect 47298 28428 47362 34572
rect -41168 22128 -41104 28272
rect -34849 22128 -34785 28272
rect -28530 22128 -28466 28272
rect -22211 22128 -22147 28272
rect -15892 22128 -15828 28272
rect -9573 22128 -9509 28272
rect -3254 22128 -3190 28272
rect 3065 22128 3129 28272
rect 9384 22128 9448 28272
rect 15703 22128 15767 28272
rect 22022 22128 22086 28272
rect 28341 22128 28405 28272
rect 34660 22128 34724 28272
rect 40979 22128 41043 28272
rect 47298 22128 47362 28272
rect -41168 15828 -41104 21972
rect -34849 15828 -34785 21972
rect -28530 15828 -28466 21972
rect -22211 15828 -22147 21972
rect -15892 15828 -15828 21972
rect -9573 15828 -9509 21972
rect -3254 15828 -3190 21972
rect 3065 15828 3129 21972
rect 9384 15828 9448 21972
rect 15703 15828 15767 21972
rect 22022 15828 22086 21972
rect 28341 15828 28405 21972
rect 34660 15828 34724 21972
rect 40979 15828 41043 21972
rect 47298 15828 47362 21972
rect -41168 9528 -41104 15672
rect -34849 9528 -34785 15672
rect -28530 9528 -28466 15672
rect -22211 9528 -22147 15672
rect -15892 9528 -15828 15672
rect -9573 9528 -9509 15672
rect -3254 9528 -3190 15672
rect 3065 9528 3129 15672
rect 9384 9528 9448 15672
rect 15703 9528 15767 15672
rect 22022 9528 22086 15672
rect 28341 9528 28405 15672
rect 34660 9528 34724 15672
rect 40979 9528 41043 15672
rect 47298 9528 47362 15672
rect -41168 3228 -41104 9372
rect -34849 3228 -34785 9372
rect -28530 3228 -28466 9372
rect -22211 3228 -22147 9372
rect -15892 3228 -15828 9372
rect -9573 3228 -9509 9372
rect -3254 3228 -3190 9372
rect 3065 3228 3129 9372
rect 9384 3228 9448 9372
rect 15703 3228 15767 9372
rect 22022 3228 22086 9372
rect 28341 3228 28405 9372
rect 34660 3228 34724 9372
rect 40979 3228 41043 9372
rect 47298 3228 47362 9372
rect -41168 -3072 -41104 3072
rect -34849 -3072 -34785 3072
rect -28530 -3072 -28466 3072
rect -22211 -3072 -22147 3072
rect -15892 -3072 -15828 3072
rect -9573 -3072 -9509 3072
rect -3254 -3072 -3190 3072
rect 3065 -3072 3129 3072
rect 9384 -3072 9448 3072
rect 15703 -3072 15767 3072
rect 22022 -3072 22086 3072
rect 28341 -3072 28405 3072
rect 34660 -3072 34724 3072
rect 40979 -3072 41043 3072
rect 47298 -3072 47362 3072
rect -41168 -9372 -41104 -3228
rect -34849 -9372 -34785 -3228
rect -28530 -9372 -28466 -3228
rect -22211 -9372 -22147 -3228
rect -15892 -9372 -15828 -3228
rect -9573 -9372 -9509 -3228
rect -3254 -9372 -3190 -3228
rect 3065 -9372 3129 -3228
rect 9384 -9372 9448 -3228
rect 15703 -9372 15767 -3228
rect 22022 -9372 22086 -3228
rect 28341 -9372 28405 -3228
rect 34660 -9372 34724 -3228
rect 40979 -9372 41043 -3228
rect 47298 -9372 47362 -3228
rect -41168 -15672 -41104 -9528
rect -34849 -15672 -34785 -9528
rect -28530 -15672 -28466 -9528
rect -22211 -15672 -22147 -9528
rect -15892 -15672 -15828 -9528
rect -9573 -15672 -9509 -9528
rect -3254 -15672 -3190 -9528
rect 3065 -15672 3129 -9528
rect 9384 -15672 9448 -9528
rect 15703 -15672 15767 -9528
rect 22022 -15672 22086 -9528
rect 28341 -15672 28405 -9528
rect 34660 -15672 34724 -9528
rect 40979 -15672 41043 -9528
rect 47298 -15672 47362 -9528
rect -41168 -21972 -41104 -15828
rect -34849 -21972 -34785 -15828
rect -28530 -21972 -28466 -15828
rect -22211 -21972 -22147 -15828
rect -15892 -21972 -15828 -15828
rect -9573 -21972 -9509 -15828
rect -3254 -21972 -3190 -15828
rect 3065 -21972 3129 -15828
rect 9384 -21972 9448 -15828
rect 15703 -21972 15767 -15828
rect 22022 -21972 22086 -15828
rect 28341 -21972 28405 -15828
rect 34660 -21972 34724 -15828
rect 40979 -21972 41043 -15828
rect 47298 -21972 47362 -15828
rect -41168 -28272 -41104 -22128
rect -34849 -28272 -34785 -22128
rect -28530 -28272 -28466 -22128
rect -22211 -28272 -22147 -22128
rect -15892 -28272 -15828 -22128
rect -9573 -28272 -9509 -22128
rect -3254 -28272 -3190 -22128
rect 3065 -28272 3129 -22128
rect 9384 -28272 9448 -22128
rect 15703 -28272 15767 -22128
rect 22022 -28272 22086 -22128
rect 28341 -28272 28405 -22128
rect 34660 -28272 34724 -22128
rect 40979 -28272 41043 -22128
rect 47298 -28272 47362 -22128
rect -41168 -34572 -41104 -28428
rect -34849 -34572 -34785 -28428
rect -28530 -34572 -28466 -28428
rect -22211 -34572 -22147 -28428
rect -15892 -34572 -15828 -28428
rect -9573 -34572 -9509 -28428
rect -3254 -34572 -3190 -28428
rect 3065 -34572 3129 -28428
rect 9384 -34572 9448 -28428
rect 15703 -34572 15767 -28428
rect 22022 -34572 22086 -28428
rect 28341 -34572 28405 -28428
rect 34660 -34572 34724 -28428
rect 40979 -34572 41043 -28428
rect 47298 -34572 47362 -28428
rect -41168 -40872 -41104 -34728
rect -34849 -40872 -34785 -34728
rect -28530 -40872 -28466 -34728
rect -22211 -40872 -22147 -34728
rect -15892 -40872 -15828 -34728
rect -9573 -40872 -9509 -34728
rect -3254 -40872 -3190 -34728
rect 3065 -40872 3129 -34728
rect 9384 -40872 9448 -34728
rect 15703 -40872 15767 -34728
rect 22022 -40872 22086 -34728
rect 28341 -40872 28405 -34728
rect 34660 -40872 34724 -34728
rect 40979 -40872 41043 -34728
rect 47298 -40872 47362 -34728
rect -41168 -47172 -41104 -41028
rect -34849 -47172 -34785 -41028
rect -28530 -47172 -28466 -41028
rect -22211 -47172 -22147 -41028
rect -15892 -47172 -15828 -41028
rect -9573 -47172 -9509 -41028
rect -3254 -47172 -3190 -41028
rect 3065 -47172 3129 -41028
rect 9384 -47172 9448 -41028
rect 15703 -47172 15767 -41028
rect 22022 -47172 22086 -41028
rect 28341 -47172 28405 -41028
rect 34660 -47172 34724 -41028
rect 40979 -47172 41043 -41028
rect 47298 -47172 47362 -41028
<< mimcap >>
rect -47283 47060 -41283 47100
rect -47283 41140 -47243 47060
rect -41323 41140 -41283 47060
rect -47283 41100 -41283 41140
rect -40964 47060 -34964 47100
rect -40964 41140 -40924 47060
rect -35004 41140 -34964 47060
rect -40964 41100 -34964 41140
rect -34645 47060 -28645 47100
rect -34645 41140 -34605 47060
rect -28685 41140 -28645 47060
rect -34645 41100 -28645 41140
rect -28326 47060 -22326 47100
rect -28326 41140 -28286 47060
rect -22366 41140 -22326 47060
rect -28326 41100 -22326 41140
rect -22007 47060 -16007 47100
rect -22007 41140 -21967 47060
rect -16047 41140 -16007 47060
rect -22007 41100 -16007 41140
rect -15688 47060 -9688 47100
rect -15688 41140 -15648 47060
rect -9728 41140 -9688 47060
rect -15688 41100 -9688 41140
rect -9369 47060 -3369 47100
rect -9369 41140 -9329 47060
rect -3409 41140 -3369 47060
rect -9369 41100 -3369 41140
rect -3050 47060 2950 47100
rect -3050 41140 -3010 47060
rect 2910 41140 2950 47060
rect -3050 41100 2950 41140
rect 3269 47060 9269 47100
rect 3269 41140 3309 47060
rect 9229 41140 9269 47060
rect 3269 41100 9269 41140
rect 9588 47060 15588 47100
rect 9588 41140 9628 47060
rect 15548 41140 15588 47060
rect 9588 41100 15588 41140
rect 15907 47060 21907 47100
rect 15907 41140 15947 47060
rect 21867 41140 21907 47060
rect 15907 41100 21907 41140
rect 22226 47060 28226 47100
rect 22226 41140 22266 47060
rect 28186 41140 28226 47060
rect 22226 41100 28226 41140
rect 28545 47060 34545 47100
rect 28545 41140 28585 47060
rect 34505 41140 34545 47060
rect 28545 41100 34545 41140
rect 34864 47060 40864 47100
rect 34864 41140 34904 47060
rect 40824 41140 40864 47060
rect 34864 41100 40864 41140
rect 41183 47060 47183 47100
rect 41183 41140 41223 47060
rect 47143 41140 47183 47060
rect 41183 41100 47183 41140
rect -47283 40760 -41283 40800
rect -47283 34840 -47243 40760
rect -41323 34840 -41283 40760
rect -47283 34800 -41283 34840
rect -40964 40760 -34964 40800
rect -40964 34840 -40924 40760
rect -35004 34840 -34964 40760
rect -40964 34800 -34964 34840
rect -34645 40760 -28645 40800
rect -34645 34840 -34605 40760
rect -28685 34840 -28645 40760
rect -34645 34800 -28645 34840
rect -28326 40760 -22326 40800
rect -28326 34840 -28286 40760
rect -22366 34840 -22326 40760
rect -28326 34800 -22326 34840
rect -22007 40760 -16007 40800
rect -22007 34840 -21967 40760
rect -16047 34840 -16007 40760
rect -22007 34800 -16007 34840
rect -15688 40760 -9688 40800
rect -15688 34840 -15648 40760
rect -9728 34840 -9688 40760
rect -15688 34800 -9688 34840
rect -9369 40760 -3369 40800
rect -9369 34840 -9329 40760
rect -3409 34840 -3369 40760
rect -9369 34800 -3369 34840
rect -3050 40760 2950 40800
rect -3050 34840 -3010 40760
rect 2910 34840 2950 40760
rect -3050 34800 2950 34840
rect 3269 40760 9269 40800
rect 3269 34840 3309 40760
rect 9229 34840 9269 40760
rect 3269 34800 9269 34840
rect 9588 40760 15588 40800
rect 9588 34840 9628 40760
rect 15548 34840 15588 40760
rect 9588 34800 15588 34840
rect 15907 40760 21907 40800
rect 15907 34840 15947 40760
rect 21867 34840 21907 40760
rect 15907 34800 21907 34840
rect 22226 40760 28226 40800
rect 22226 34840 22266 40760
rect 28186 34840 28226 40760
rect 22226 34800 28226 34840
rect 28545 40760 34545 40800
rect 28545 34840 28585 40760
rect 34505 34840 34545 40760
rect 28545 34800 34545 34840
rect 34864 40760 40864 40800
rect 34864 34840 34904 40760
rect 40824 34840 40864 40760
rect 34864 34800 40864 34840
rect 41183 40760 47183 40800
rect 41183 34840 41223 40760
rect 47143 34840 47183 40760
rect 41183 34800 47183 34840
rect -47283 34460 -41283 34500
rect -47283 28540 -47243 34460
rect -41323 28540 -41283 34460
rect -47283 28500 -41283 28540
rect -40964 34460 -34964 34500
rect -40964 28540 -40924 34460
rect -35004 28540 -34964 34460
rect -40964 28500 -34964 28540
rect -34645 34460 -28645 34500
rect -34645 28540 -34605 34460
rect -28685 28540 -28645 34460
rect -34645 28500 -28645 28540
rect -28326 34460 -22326 34500
rect -28326 28540 -28286 34460
rect -22366 28540 -22326 34460
rect -28326 28500 -22326 28540
rect -22007 34460 -16007 34500
rect -22007 28540 -21967 34460
rect -16047 28540 -16007 34460
rect -22007 28500 -16007 28540
rect -15688 34460 -9688 34500
rect -15688 28540 -15648 34460
rect -9728 28540 -9688 34460
rect -15688 28500 -9688 28540
rect -9369 34460 -3369 34500
rect -9369 28540 -9329 34460
rect -3409 28540 -3369 34460
rect -9369 28500 -3369 28540
rect -3050 34460 2950 34500
rect -3050 28540 -3010 34460
rect 2910 28540 2950 34460
rect -3050 28500 2950 28540
rect 3269 34460 9269 34500
rect 3269 28540 3309 34460
rect 9229 28540 9269 34460
rect 3269 28500 9269 28540
rect 9588 34460 15588 34500
rect 9588 28540 9628 34460
rect 15548 28540 15588 34460
rect 9588 28500 15588 28540
rect 15907 34460 21907 34500
rect 15907 28540 15947 34460
rect 21867 28540 21907 34460
rect 15907 28500 21907 28540
rect 22226 34460 28226 34500
rect 22226 28540 22266 34460
rect 28186 28540 28226 34460
rect 22226 28500 28226 28540
rect 28545 34460 34545 34500
rect 28545 28540 28585 34460
rect 34505 28540 34545 34460
rect 28545 28500 34545 28540
rect 34864 34460 40864 34500
rect 34864 28540 34904 34460
rect 40824 28540 40864 34460
rect 34864 28500 40864 28540
rect 41183 34460 47183 34500
rect 41183 28540 41223 34460
rect 47143 28540 47183 34460
rect 41183 28500 47183 28540
rect -47283 28160 -41283 28200
rect -47283 22240 -47243 28160
rect -41323 22240 -41283 28160
rect -47283 22200 -41283 22240
rect -40964 28160 -34964 28200
rect -40964 22240 -40924 28160
rect -35004 22240 -34964 28160
rect -40964 22200 -34964 22240
rect -34645 28160 -28645 28200
rect -34645 22240 -34605 28160
rect -28685 22240 -28645 28160
rect -34645 22200 -28645 22240
rect -28326 28160 -22326 28200
rect -28326 22240 -28286 28160
rect -22366 22240 -22326 28160
rect -28326 22200 -22326 22240
rect -22007 28160 -16007 28200
rect -22007 22240 -21967 28160
rect -16047 22240 -16007 28160
rect -22007 22200 -16007 22240
rect -15688 28160 -9688 28200
rect -15688 22240 -15648 28160
rect -9728 22240 -9688 28160
rect -15688 22200 -9688 22240
rect -9369 28160 -3369 28200
rect -9369 22240 -9329 28160
rect -3409 22240 -3369 28160
rect -9369 22200 -3369 22240
rect -3050 28160 2950 28200
rect -3050 22240 -3010 28160
rect 2910 22240 2950 28160
rect -3050 22200 2950 22240
rect 3269 28160 9269 28200
rect 3269 22240 3309 28160
rect 9229 22240 9269 28160
rect 3269 22200 9269 22240
rect 9588 28160 15588 28200
rect 9588 22240 9628 28160
rect 15548 22240 15588 28160
rect 9588 22200 15588 22240
rect 15907 28160 21907 28200
rect 15907 22240 15947 28160
rect 21867 22240 21907 28160
rect 15907 22200 21907 22240
rect 22226 28160 28226 28200
rect 22226 22240 22266 28160
rect 28186 22240 28226 28160
rect 22226 22200 28226 22240
rect 28545 28160 34545 28200
rect 28545 22240 28585 28160
rect 34505 22240 34545 28160
rect 28545 22200 34545 22240
rect 34864 28160 40864 28200
rect 34864 22240 34904 28160
rect 40824 22240 40864 28160
rect 34864 22200 40864 22240
rect 41183 28160 47183 28200
rect 41183 22240 41223 28160
rect 47143 22240 47183 28160
rect 41183 22200 47183 22240
rect -47283 21860 -41283 21900
rect -47283 15940 -47243 21860
rect -41323 15940 -41283 21860
rect -47283 15900 -41283 15940
rect -40964 21860 -34964 21900
rect -40964 15940 -40924 21860
rect -35004 15940 -34964 21860
rect -40964 15900 -34964 15940
rect -34645 21860 -28645 21900
rect -34645 15940 -34605 21860
rect -28685 15940 -28645 21860
rect -34645 15900 -28645 15940
rect -28326 21860 -22326 21900
rect -28326 15940 -28286 21860
rect -22366 15940 -22326 21860
rect -28326 15900 -22326 15940
rect -22007 21860 -16007 21900
rect -22007 15940 -21967 21860
rect -16047 15940 -16007 21860
rect -22007 15900 -16007 15940
rect -15688 21860 -9688 21900
rect -15688 15940 -15648 21860
rect -9728 15940 -9688 21860
rect -15688 15900 -9688 15940
rect -9369 21860 -3369 21900
rect -9369 15940 -9329 21860
rect -3409 15940 -3369 21860
rect -9369 15900 -3369 15940
rect -3050 21860 2950 21900
rect -3050 15940 -3010 21860
rect 2910 15940 2950 21860
rect -3050 15900 2950 15940
rect 3269 21860 9269 21900
rect 3269 15940 3309 21860
rect 9229 15940 9269 21860
rect 3269 15900 9269 15940
rect 9588 21860 15588 21900
rect 9588 15940 9628 21860
rect 15548 15940 15588 21860
rect 9588 15900 15588 15940
rect 15907 21860 21907 21900
rect 15907 15940 15947 21860
rect 21867 15940 21907 21860
rect 15907 15900 21907 15940
rect 22226 21860 28226 21900
rect 22226 15940 22266 21860
rect 28186 15940 28226 21860
rect 22226 15900 28226 15940
rect 28545 21860 34545 21900
rect 28545 15940 28585 21860
rect 34505 15940 34545 21860
rect 28545 15900 34545 15940
rect 34864 21860 40864 21900
rect 34864 15940 34904 21860
rect 40824 15940 40864 21860
rect 34864 15900 40864 15940
rect 41183 21860 47183 21900
rect 41183 15940 41223 21860
rect 47143 15940 47183 21860
rect 41183 15900 47183 15940
rect -47283 15560 -41283 15600
rect -47283 9640 -47243 15560
rect -41323 9640 -41283 15560
rect -47283 9600 -41283 9640
rect -40964 15560 -34964 15600
rect -40964 9640 -40924 15560
rect -35004 9640 -34964 15560
rect -40964 9600 -34964 9640
rect -34645 15560 -28645 15600
rect -34645 9640 -34605 15560
rect -28685 9640 -28645 15560
rect -34645 9600 -28645 9640
rect -28326 15560 -22326 15600
rect -28326 9640 -28286 15560
rect -22366 9640 -22326 15560
rect -28326 9600 -22326 9640
rect -22007 15560 -16007 15600
rect -22007 9640 -21967 15560
rect -16047 9640 -16007 15560
rect -22007 9600 -16007 9640
rect -15688 15560 -9688 15600
rect -15688 9640 -15648 15560
rect -9728 9640 -9688 15560
rect -15688 9600 -9688 9640
rect -9369 15560 -3369 15600
rect -9369 9640 -9329 15560
rect -3409 9640 -3369 15560
rect -9369 9600 -3369 9640
rect -3050 15560 2950 15600
rect -3050 9640 -3010 15560
rect 2910 9640 2950 15560
rect -3050 9600 2950 9640
rect 3269 15560 9269 15600
rect 3269 9640 3309 15560
rect 9229 9640 9269 15560
rect 3269 9600 9269 9640
rect 9588 15560 15588 15600
rect 9588 9640 9628 15560
rect 15548 9640 15588 15560
rect 9588 9600 15588 9640
rect 15907 15560 21907 15600
rect 15907 9640 15947 15560
rect 21867 9640 21907 15560
rect 15907 9600 21907 9640
rect 22226 15560 28226 15600
rect 22226 9640 22266 15560
rect 28186 9640 28226 15560
rect 22226 9600 28226 9640
rect 28545 15560 34545 15600
rect 28545 9640 28585 15560
rect 34505 9640 34545 15560
rect 28545 9600 34545 9640
rect 34864 15560 40864 15600
rect 34864 9640 34904 15560
rect 40824 9640 40864 15560
rect 34864 9600 40864 9640
rect 41183 15560 47183 15600
rect 41183 9640 41223 15560
rect 47143 9640 47183 15560
rect 41183 9600 47183 9640
rect -47283 9260 -41283 9300
rect -47283 3340 -47243 9260
rect -41323 3340 -41283 9260
rect -47283 3300 -41283 3340
rect -40964 9260 -34964 9300
rect -40964 3340 -40924 9260
rect -35004 3340 -34964 9260
rect -40964 3300 -34964 3340
rect -34645 9260 -28645 9300
rect -34645 3340 -34605 9260
rect -28685 3340 -28645 9260
rect -34645 3300 -28645 3340
rect -28326 9260 -22326 9300
rect -28326 3340 -28286 9260
rect -22366 3340 -22326 9260
rect -28326 3300 -22326 3340
rect -22007 9260 -16007 9300
rect -22007 3340 -21967 9260
rect -16047 3340 -16007 9260
rect -22007 3300 -16007 3340
rect -15688 9260 -9688 9300
rect -15688 3340 -15648 9260
rect -9728 3340 -9688 9260
rect -15688 3300 -9688 3340
rect -9369 9260 -3369 9300
rect -9369 3340 -9329 9260
rect -3409 3340 -3369 9260
rect -9369 3300 -3369 3340
rect -3050 9260 2950 9300
rect -3050 3340 -3010 9260
rect 2910 3340 2950 9260
rect -3050 3300 2950 3340
rect 3269 9260 9269 9300
rect 3269 3340 3309 9260
rect 9229 3340 9269 9260
rect 3269 3300 9269 3340
rect 9588 9260 15588 9300
rect 9588 3340 9628 9260
rect 15548 3340 15588 9260
rect 9588 3300 15588 3340
rect 15907 9260 21907 9300
rect 15907 3340 15947 9260
rect 21867 3340 21907 9260
rect 15907 3300 21907 3340
rect 22226 9260 28226 9300
rect 22226 3340 22266 9260
rect 28186 3340 28226 9260
rect 22226 3300 28226 3340
rect 28545 9260 34545 9300
rect 28545 3340 28585 9260
rect 34505 3340 34545 9260
rect 28545 3300 34545 3340
rect 34864 9260 40864 9300
rect 34864 3340 34904 9260
rect 40824 3340 40864 9260
rect 34864 3300 40864 3340
rect 41183 9260 47183 9300
rect 41183 3340 41223 9260
rect 47143 3340 47183 9260
rect 41183 3300 47183 3340
rect -47283 2960 -41283 3000
rect -47283 -2960 -47243 2960
rect -41323 -2960 -41283 2960
rect -47283 -3000 -41283 -2960
rect -40964 2960 -34964 3000
rect -40964 -2960 -40924 2960
rect -35004 -2960 -34964 2960
rect -40964 -3000 -34964 -2960
rect -34645 2960 -28645 3000
rect -34645 -2960 -34605 2960
rect -28685 -2960 -28645 2960
rect -34645 -3000 -28645 -2960
rect -28326 2960 -22326 3000
rect -28326 -2960 -28286 2960
rect -22366 -2960 -22326 2960
rect -28326 -3000 -22326 -2960
rect -22007 2960 -16007 3000
rect -22007 -2960 -21967 2960
rect -16047 -2960 -16007 2960
rect -22007 -3000 -16007 -2960
rect -15688 2960 -9688 3000
rect -15688 -2960 -15648 2960
rect -9728 -2960 -9688 2960
rect -15688 -3000 -9688 -2960
rect -9369 2960 -3369 3000
rect -9369 -2960 -9329 2960
rect -3409 -2960 -3369 2960
rect -9369 -3000 -3369 -2960
rect -3050 2960 2950 3000
rect -3050 -2960 -3010 2960
rect 2910 -2960 2950 2960
rect -3050 -3000 2950 -2960
rect 3269 2960 9269 3000
rect 3269 -2960 3309 2960
rect 9229 -2960 9269 2960
rect 3269 -3000 9269 -2960
rect 9588 2960 15588 3000
rect 9588 -2960 9628 2960
rect 15548 -2960 15588 2960
rect 9588 -3000 15588 -2960
rect 15907 2960 21907 3000
rect 15907 -2960 15947 2960
rect 21867 -2960 21907 2960
rect 15907 -3000 21907 -2960
rect 22226 2960 28226 3000
rect 22226 -2960 22266 2960
rect 28186 -2960 28226 2960
rect 22226 -3000 28226 -2960
rect 28545 2960 34545 3000
rect 28545 -2960 28585 2960
rect 34505 -2960 34545 2960
rect 28545 -3000 34545 -2960
rect 34864 2960 40864 3000
rect 34864 -2960 34904 2960
rect 40824 -2960 40864 2960
rect 34864 -3000 40864 -2960
rect 41183 2960 47183 3000
rect 41183 -2960 41223 2960
rect 47143 -2960 47183 2960
rect 41183 -3000 47183 -2960
rect -47283 -3340 -41283 -3300
rect -47283 -9260 -47243 -3340
rect -41323 -9260 -41283 -3340
rect -47283 -9300 -41283 -9260
rect -40964 -3340 -34964 -3300
rect -40964 -9260 -40924 -3340
rect -35004 -9260 -34964 -3340
rect -40964 -9300 -34964 -9260
rect -34645 -3340 -28645 -3300
rect -34645 -9260 -34605 -3340
rect -28685 -9260 -28645 -3340
rect -34645 -9300 -28645 -9260
rect -28326 -3340 -22326 -3300
rect -28326 -9260 -28286 -3340
rect -22366 -9260 -22326 -3340
rect -28326 -9300 -22326 -9260
rect -22007 -3340 -16007 -3300
rect -22007 -9260 -21967 -3340
rect -16047 -9260 -16007 -3340
rect -22007 -9300 -16007 -9260
rect -15688 -3340 -9688 -3300
rect -15688 -9260 -15648 -3340
rect -9728 -9260 -9688 -3340
rect -15688 -9300 -9688 -9260
rect -9369 -3340 -3369 -3300
rect -9369 -9260 -9329 -3340
rect -3409 -9260 -3369 -3340
rect -9369 -9300 -3369 -9260
rect -3050 -3340 2950 -3300
rect -3050 -9260 -3010 -3340
rect 2910 -9260 2950 -3340
rect -3050 -9300 2950 -9260
rect 3269 -3340 9269 -3300
rect 3269 -9260 3309 -3340
rect 9229 -9260 9269 -3340
rect 3269 -9300 9269 -9260
rect 9588 -3340 15588 -3300
rect 9588 -9260 9628 -3340
rect 15548 -9260 15588 -3340
rect 9588 -9300 15588 -9260
rect 15907 -3340 21907 -3300
rect 15907 -9260 15947 -3340
rect 21867 -9260 21907 -3340
rect 15907 -9300 21907 -9260
rect 22226 -3340 28226 -3300
rect 22226 -9260 22266 -3340
rect 28186 -9260 28226 -3340
rect 22226 -9300 28226 -9260
rect 28545 -3340 34545 -3300
rect 28545 -9260 28585 -3340
rect 34505 -9260 34545 -3340
rect 28545 -9300 34545 -9260
rect 34864 -3340 40864 -3300
rect 34864 -9260 34904 -3340
rect 40824 -9260 40864 -3340
rect 34864 -9300 40864 -9260
rect 41183 -3340 47183 -3300
rect 41183 -9260 41223 -3340
rect 47143 -9260 47183 -3340
rect 41183 -9300 47183 -9260
rect -47283 -9640 -41283 -9600
rect -47283 -15560 -47243 -9640
rect -41323 -15560 -41283 -9640
rect -47283 -15600 -41283 -15560
rect -40964 -9640 -34964 -9600
rect -40964 -15560 -40924 -9640
rect -35004 -15560 -34964 -9640
rect -40964 -15600 -34964 -15560
rect -34645 -9640 -28645 -9600
rect -34645 -15560 -34605 -9640
rect -28685 -15560 -28645 -9640
rect -34645 -15600 -28645 -15560
rect -28326 -9640 -22326 -9600
rect -28326 -15560 -28286 -9640
rect -22366 -15560 -22326 -9640
rect -28326 -15600 -22326 -15560
rect -22007 -9640 -16007 -9600
rect -22007 -15560 -21967 -9640
rect -16047 -15560 -16007 -9640
rect -22007 -15600 -16007 -15560
rect -15688 -9640 -9688 -9600
rect -15688 -15560 -15648 -9640
rect -9728 -15560 -9688 -9640
rect -15688 -15600 -9688 -15560
rect -9369 -9640 -3369 -9600
rect -9369 -15560 -9329 -9640
rect -3409 -15560 -3369 -9640
rect -9369 -15600 -3369 -15560
rect -3050 -9640 2950 -9600
rect -3050 -15560 -3010 -9640
rect 2910 -15560 2950 -9640
rect -3050 -15600 2950 -15560
rect 3269 -9640 9269 -9600
rect 3269 -15560 3309 -9640
rect 9229 -15560 9269 -9640
rect 3269 -15600 9269 -15560
rect 9588 -9640 15588 -9600
rect 9588 -15560 9628 -9640
rect 15548 -15560 15588 -9640
rect 9588 -15600 15588 -15560
rect 15907 -9640 21907 -9600
rect 15907 -15560 15947 -9640
rect 21867 -15560 21907 -9640
rect 15907 -15600 21907 -15560
rect 22226 -9640 28226 -9600
rect 22226 -15560 22266 -9640
rect 28186 -15560 28226 -9640
rect 22226 -15600 28226 -15560
rect 28545 -9640 34545 -9600
rect 28545 -15560 28585 -9640
rect 34505 -15560 34545 -9640
rect 28545 -15600 34545 -15560
rect 34864 -9640 40864 -9600
rect 34864 -15560 34904 -9640
rect 40824 -15560 40864 -9640
rect 34864 -15600 40864 -15560
rect 41183 -9640 47183 -9600
rect 41183 -15560 41223 -9640
rect 47143 -15560 47183 -9640
rect 41183 -15600 47183 -15560
rect -47283 -15940 -41283 -15900
rect -47283 -21860 -47243 -15940
rect -41323 -21860 -41283 -15940
rect -47283 -21900 -41283 -21860
rect -40964 -15940 -34964 -15900
rect -40964 -21860 -40924 -15940
rect -35004 -21860 -34964 -15940
rect -40964 -21900 -34964 -21860
rect -34645 -15940 -28645 -15900
rect -34645 -21860 -34605 -15940
rect -28685 -21860 -28645 -15940
rect -34645 -21900 -28645 -21860
rect -28326 -15940 -22326 -15900
rect -28326 -21860 -28286 -15940
rect -22366 -21860 -22326 -15940
rect -28326 -21900 -22326 -21860
rect -22007 -15940 -16007 -15900
rect -22007 -21860 -21967 -15940
rect -16047 -21860 -16007 -15940
rect -22007 -21900 -16007 -21860
rect -15688 -15940 -9688 -15900
rect -15688 -21860 -15648 -15940
rect -9728 -21860 -9688 -15940
rect -15688 -21900 -9688 -21860
rect -9369 -15940 -3369 -15900
rect -9369 -21860 -9329 -15940
rect -3409 -21860 -3369 -15940
rect -9369 -21900 -3369 -21860
rect -3050 -15940 2950 -15900
rect -3050 -21860 -3010 -15940
rect 2910 -21860 2950 -15940
rect -3050 -21900 2950 -21860
rect 3269 -15940 9269 -15900
rect 3269 -21860 3309 -15940
rect 9229 -21860 9269 -15940
rect 3269 -21900 9269 -21860
rect 9588 -15940 15588 -15900
rect 9588 -21860 9628 -15940
rect 15548 -21860 15588 -15940
rect 9588 -21900 15588 -21860
rect 15907 -15940 21907 -15900
rect 15907 -21860 15947 -15940
rect 21867 -21860 21907 -15940
rect 15907 -21900 21907 -21860
rect 22226 -15940 28226 -15900
rect 22226 -21860 22266 -15940
rect 28186 -21860 28226 -15940
rect 22226 -21900 28226 -21860
rect 28545 -15940 34545 -15900
rect 28545 -21860 28585 -15940
rect 34505 -21860 34545 -15940
rect 28545 -21900 34545 -21860
rect 34864 -15940 40864 -15900
rect 34864 -21860 34904 -15940
rect 40824 -21860 40864 -15940
rect 34864 -21900 40864 -21860
rect 41183 -15940 47183 -15900
rect 41183 -21860 41223 -15940
rect 47143 -21860 47183 -15940
rect 41183 -21900 47183 -21860
rect -47283 -22240 -41283 -22200
rect -47283 -28160 -47243 -22240
rect -41323 -28160 -41283 -22240
rect -47283 -28200 -41283 -28160
rect -40964 -22240 -34964 -22200
rect -40964 -28160 -40924 -22240
rect -35004 -28160 -34964 -22240
rect -40964 -28200 -34964 -28160
rect -34645 -22240 -28645 -22200
rect -34645 -28160 -34605 -22240
rect -28685 -28160 -28645 -22240
rect -34645 -28200 -28645 -28160
rect -28326 -22240 -22326 -22200
rect -28326 -28160 -28286 -22240
rect -22366 -28160 -22326 -22240
rect -28326 -28200 -22326 -28160
rect -22007 -22240 -16007 -22200
rect -22007 -28160 -21967 -22240
rect -16047 -28160 -16007 -22240
rect -22007 -28200 -16007 -28160
rect -15688 -22240 -9688 -22200
rect -15688 -28160 -15648 -22240
rect -9728 -28160 -9688 -22240
rect -15688 -28200 -9688 -28160
rect -9369 -22240 -3369 -22200
rect -9369 -28160 -9329 -22240
rect -3409 -28160 -3369 -22240
rect -9369 -28200 -3369 -28160
rect -3050 -22240 2950 -22200
rect -3050 -28160 -3010 -22240
rect 2910 -28160 2950 -22240
rect -3050 -28200 2950 -28160
rect 3269 -22240 9269 -22200
rect 3269 -28160 3309 -22240
rect 9229 -28160 9269 -22240
rect 3269 -28200 9269 -28160
rect 9588 -22240 15588 -22200
rect 9588 -28160 9628 -22240
rect 15548 -28160 15588 -22240
rect 9588 -28200 15588 -28160
rect 15907 -22240 21907 -22200
rect 15907 -28160 15947 -22240
rect 21867 -28160 21907 -22240
rect 15907 -28200 21907 -28160
rect 22226 -22240 28226 -22200
rect 22226 -28160 22266 -22240
rect 28186 -28160 28226 -22240
rect 22226 -28200 28226 -28160
rect 28545 -22240 34545 -22200
rect 28545 -28160 28585 -22240
rect 34505 -28160 34545 -22240
rect 28545 -28200 34545 -28160
rect 34864 -22240 40864 -22200
rect 34864 -28160 34904 -22240
rect 40824 -28160 40864 -22240
rect 34864 -28200 40864 -28160
rect 41183 -22240 47183 -22200
rect 41183 -28160 41223 -22240
rect 47143 -28160 47183 -22240
rect 41183 -28200 47183 -28160
rect -47283 -28540 -41283 -28500
rect -47283 -34460 -47243 -28540
rect -41323 -34460 -41283 -28540
rect -47283 -34500 -41283 -34460
rect -40964 -28540 -34964 -28500
rect -40964 -34460 -40924 -28540
rect -35004 -34460 -34964 -28540
rect -40964 -34500 -34964 -34460
rect -34645 -28540 -28645 -28500
rect -34645 -34460 -34605 -28540
rect -28685 -34460 -28645 -28540
rect -34645 -34500 -28645 -34460
rect -28326 -28540 -22326 -28500
rect -28326 -34460 -28286 -28540
rect -22366 -34460 -22326 -28540
rect -28326 -34500 -22326 -34460
rect -22007 -28540 -16007 -28500
rect -22007 -34460 -21967 -28540
rect -16047 -34460 -16007 -28540
rect -22007 -34500 -16007 -34460
rect -15688 -28540 -9688 -28500
rect -15688 -34460 -15648 -28540
rect -9728 -34460 -9688 -28540
rect -15688 -34500 -9688 -34460
rect -9369 -28540 -3369 -28500
rect -9369 -34460 -9329 -28540
rect -3409 -34460 -3369 -28540
rect -9369 -34500 -3369 -34460
rect -3050 -28540 2950 -28500
rect -3050 -34460 -3010 -28540
rect 2910 -34460 2950 -28540
rect -3050 -34500 2950 -34460
rect 3269 -28540 9269 -28500
rect 3269 -34460 3309 -28540
rect 9229 -34460 9269 -28540
rect 3269 -34500 9269 -34460
rect 9588 -28540 15588 -28500
rect 9588 -34460 9628 -28540
rect 15548 -34460 15588 -28540
rect 9588 -34500 15588 -34460
rect 15907 -28540 21907 -28500
rect 15907 -34460 15947 -28540
rect 21867 -34460 21907 -28540
rect 15907 -34500 21907 -34460
rect 22226 -28540 28226 -28500
rect 22226 -34460 22266 -28540
rect 28186 -34460 28226 -28540
rect 22226 -34500 28226 -34460
rect 28545 -28540 34545 -28500
rect 28545 -34460 28585 -28540
rect 34505 -34460 34545 -28540
rect 28545 -34500 34545 -34460
rect 34864 -28540 40864 -28500
rect 34864 -34460 34904 -28540
rect 40824 -34460 40864 -28540
rect 34864 -34500 40864 -34460
rect 41183 -28540 47183 -28500
rect 41183 -34460 41223 -28540
rect 47143 -34460 47183 -28540
rect 41183 -34500 47183 -34460
rect -47283 -34840 -41283 -34800
rect -47283 -40760 -47243 -34840
rect -41323 -40760 -41283 -34840
rect -47283 -40800 -41283 -40760
rect -40964 -34840 -34964 -34800
rect -40964 -40760 -40924 -34840
rect -35004 -40760 -34964 -34840
rect -40964 -40800 -34964 -40760
rect -34645 -34840 -28645 -34800
rect -34645 -40760 -34605 -34840
rect -28685 -40760 -28645 -34840
rect -34645 -40800 -28645 -40760
rect -28326 -34840 -22326 -34800
rect -28326 -40760 -28286 -34840
rect -22366 -40760 -22326 -34840
rect -28326 -40800 -22326 -40760
rect -22007 -34840 -16007 -34800
rect -22007 -40760 -21967 -34840
rect -16047 -40760 -16007 -34840
rect -22007 -40800 -16007 -40760
rect -15688 -34840 -9688 -34800
rect -15688 -40760 -15648 -34840
rect -9728 -40760 -9688 -34840
rect -15688 -40800 -9688 -40760
rect -9369 -34840 -3369 -34800
rect -9369 -40760 -9329 -34840
rect -3409 -40760 -3369 -34840
rect -9369 -40800 -3369 -40760
rect -3050 -34840 2950 -34800
rect -3050 -40760 -3010 -34840
rect 2910 -40760 2950 -34840
rect -3050 -40800 2950 -40760
rect 3269 -34840 9269 -34800
rect 3269 -40760 3309 -34840
rect 9229 -40760 9269 -34840
rect 3269 -40800 9269 -40760
rect 9588 -34840 15588 -34800
rect 9588 -40760 9628 -34840
rect 15548 -40760 15588 -34840
rect 9588 -40800 15588 -40760
rect 15907 -34840 21907 -34800
rect 15907 -40760 15947 -34840
rect 21867 -40760 21907 -34840
rect 15907 -40800 21907 -40760
rect 22226 -34840 28226 -34800
rect 22226 -40760 22266 -34840
rect 28186 -40760 28226 -34840
rect 22226 -40800 28226 -40760
rect 28545 -34840 34545 -34800
rect 28545 -40760 28585 -34840
rect 34505 -40760 34545 -34840
rect 28545 -40800 34545 -40760
rect 34864 -34840 40864 -34800
rect 34864 -40760 34904 -34840
rect 40824 -40760 40864 -34840
rect 34864 -40800 40864 -40760
rect 41183 -34840 47183 -34800
rect 41183 -40760 41223 -34840
rect 47143 -40760 47183 -34840
rect 41183 -40800 47183 -40760
rect -47283 -41140 -41283 -41100
rect -47283 -47060 -47243 -41140
rect -41323 -47060 -41283 -41140
rect -47283 -47100 -41283 -47060
rect -40964 -41140 -34964 -41100
rect -40964 -47060 -40924 -41140
rect -35004 -47060 -34964 -41140
rect -40964 -47100 -34964 -47060
rect -34645 -41140 -28645 -41100
rect -34645 -47060 -34605 -41140
rect -28685 -47060 -28645 -41140
rect -34645 -47100 -28645 -47060
rect -28326 -41140 -22326 -41100
rect -28326 -47060 -28286 -41140
rect -22366 -47060 -22326 -41140
rect -28326 -47100 -22326 -47060
rect -22007 -41140 -16007 -41100
rect -22007 -47060 -21967 -41140
rect -16047 -47060 -16007 -41140
rect -22007 -47100 -16007 -47060
rect -15688 -41140 -9688 -41100
rect -15688 -47060 -15648 -41140
rect -9728 -47060 -9688 -41140
rect -15688 -47100 -9688 -47060
rect -9369 -41140 -3369 -41100
rect -9369 -47060 -9329 -41140
rect -3409 -47060 -3369 -41140
rect -9369 -47100 -3369 -47060
rect -3050 -41140 2950 -41100
rect -3050 -47060 -3010 -41140
rect 2910 -47060 2950 -41140
rect -3050 -47100 2950 -47060
rect 3269 -41140 9269 -41100
rect 3269 -47060 3309 -41140
rect 9229 -47060 9269 -41140
rect 3269 -47100 9269 -47060
rect 9588 -41140 15588 -41100
rect 9588 -47060 9628 -41140
rect 15548 -47060 15588 -41140
rect 9588 -47100 15588 -47060
rect 15907 -41140 21907 -41100
rect 15907 -47060 15947 -41140
rect 21867 -47060 21907 -41140
rect 15907 -47100 21907 -47060
rect 22226 -41140 28226 -41100
rect 22226 -47060 22266 -41140
rect 28186 -47060 28226 -41140
rect 22226 -47100 28226 -47060
rect 28545 -41140 34545 -41100
rect 28545 -47060 28585 -41140
rect 34505 -47060 34545 -41140
rect 28545 -47100 34545 -47060
rect 34864 -41140 40864 -41100
rect 34864 -47060 34904 -41140
rect 40824 -47060 40864 -41140
rect 34864 -47100 40864 -47060
rect 41183 -41140 47183 -41100
rect 41183 -47060 41223 -41140
rect 47143 -47060 47183 -41140
rect 41183 -47100 47183 -47060
<< mimcapcontact >>
rect -47243 41140 -41323 47060
rect -40924 41140 -35004 47060
rect -34605 41140 -28685 47060
rect -28286 41140 -22366 47060
rect -21967 41140 -16047 47060
rect -15648 41140 -9728 47060
rect -9329 41140 -3409 47060
rect -3010 41140 2910 47060
rect 3309 41140 9229 47060
rect 9628 41140 15548 47060
rect 15947 41140 21867 47060
rect 22266 41140 28186 47060
rect 28585 41140 34505 47060
rect 34904 41140 40824 47060
rect 41223 41140 47143 47060
rect -47243 34840 -41323 40760
rect -40924 34840 -35004 40760
rect -34605 34840 -28685 40760
rect -28286 34840 -22366 40760
rect -21967 34840 -16047 40760
rect -15648 34840 -9728 40760
rect -9329 34840 -3409 40760
rect -3010 34840 2910 40760
rect 3309 34840 9229 40760
rect 9628 34840 15548 40760
rect 15947 34840 21867 40760
rect 22266 34840 28186 40760
rect 28585 34840 34505 40760
rect 34904 34840 40824 40760
rect 41223 34840 47143 40760
rect -47243 28540 -41323 34460
rect -40924 28540 -35004 34460
rect -34605 28540 -28685 34460
rect -28286 28540 -22366 34460
rect -21967 28540 -16047 34460
rect -15648 28540 -9728 34460
rect -9329 28540 -3409 34460
rect -3010 28540 2910 34460
rect 3309 28540 9229 34460
rect 9628 28540 15548 34460
rect 15947 28540 21867 34460
rect 22266 28540 28186 34460
rect 28585 28540 34505 34460
rect 34904 28540 40824 34460
rect 41223 28540 47143 34460
rect -47243 22240 -41323 28160
rect -40924 22240 -35004 28160
rect -34605 22240 -28685 28160
rect -28286 22240 -22366 28160
rect -21967 22240 -16047 28160
rect -15648 22240 -9728 28160
rect -9329 22240 -3409 28160
rect -3010 22240 2910 28160
rect 3309 22240 9229 28160
rect 9628 22240 15548 28160
rect 15947 22240 21867 28160
rect 22266 22240 28186 28160
rect 28585 22240 34505 28160
rect 34904 22240 40824 28160
rect 41223 22240 47143 28160
rect -47243 15940 -41323 21860
rect -40924 15940 -35004 21860
rect -34605 15940 -28685 21860
rect -28286 15940 -22366 21860
rect -21967 15940 -16047 21860
rect -15648 15940 -9728 21860
rect -9329 15940 -3409 21860
rect -3010 15940 2910 21860
rect 3309 15940 9229 21860
rect 9628 15940 15548 21860
rect 15947 15940 21867 21860
rect 22266 15940 28186 21860
rect 28585 15940 34505 21860
rect 34904 15940 40824 21860
rect 41223 15940 47143 21860
rect -47243 9640 -41323 15560
rect -40924 9640 -35004 15560
rect -34605 9640 -28685 15560
rect -28286 9640 -22366 15560
rect -21967 9640 -16047 15560
rect -15648 9640 -9728 15560
rect -9329 9640 -3409 15560
rect -3010 9640 2910 15560
rect 3309 9640 9229 15560
rect 9628 9640 15548 15560
rect 15947 9640 21867 15560
rect 22266 9640 28186 15560
rect 28585 9640 34505 15560
rect 34904 9640 40824 15560
rect 41223 9640 47143 15560
rect -47243 3340 -41323 9260
rect -40924 3340 -35004 9260
rect -34605 3340 -28685 9260
rect -28286 3340 -22366 9260
rect -21967 3340 -16047 9260
rect -15648 3340 -9728 9260
rect -9329 3340 -3409 9260
rect -3010 3340 2910 9260
rect 3309 3340 9229 9260
rect 9628 3340 15548 9260
rect 15947 3340 21867 9260
rect 22266 3340 28186 9260
rect 28585 3340 34505 9260
rect 34904 3340 40824 9260
rect 41223 3340 47143 9260
rect -47243 -2960 -41323 2960
rect -40924 -2960 -35004 2960
rect -34605 -2960 -28685 2960
rect -28286 -2960 -22366 2960
rect -21967 -2960 -16047 2960
rect -15648 -2960 -9728 2960
rect -9329 -2960 -3409 2960
rect -3010 -2960 2910 2960
rect 3309 -2960 9229 2960
rect 9628 -2960 15548 2960
rect 15947 -2960 21867 2960
rect 22266 -2960 28186 2960
rect 28585 -2960 34505 2960
rect 34904 -2960 40824 2960
rect 41223 -2960 47143 2960
rect -47243 -9260 -41323 -3340
rect -40924 -9260 -35004 -3340
rect -34605 -9260 -28685 -3340
rect -28286 -9260 -22366 -3340
rect -21967 -9260 -16047 -3340
rect -15648 -9260 -9728 -3340
rect -9329 -9260 -3409 -3340
rect -3010 -9260 2910 -3340
rect 3309 -9260 9229 -3340
rect 9628 -9260 15548 -3340
rect 15947 -9260 21867 -3340
rect 22266 -9260 28186 -3340
rect 28585 -9260 34505 -3340
rect 34904 -9260 40824 -3340
rect 41223 -9260 47143 -3340
rect -47243 -15560 -41323 -9640
rect -40924 -15560 -35004 -9640
rect -34605 -15560 -28685 -9640
rect -28286 -15560 -22366 -9640
rect -21967 -15560 -16047 -9640
rect -15648 -15560 -9728 -9640
rect -9329 -15560 -3409 -9640
rect -3010 -15560 2910 -9640
rect 3309 -15560 9229 -9640
rect 9628 -15560 15548 -9640
rect 15947 -15560 21867 -9640
rect 22266 -15560 28186 -9640
rect 28585 -15560 34505 -9640
rect 34904 -15560 40824 -9640
rect 41223 -15560 47143 -9640
rect -47243 -21860 -41323 -15940
rect -40924 -21860 -35004 -15940
rect -34605 -21860 -28685 -15940
rect -28286 -21860 -22366 -15940
rect -21967 -21860 -16047 -15940
rect -15648 -21860 -9728 -15940
rect -9329 -21860 -3409 -15940
rect -3010 -21860 2910 -15940
rect 3309 -21860 9229 -15940
rect 9628 -21860 15548 -15940
rect 15947 -21860 21867 -15940
rect 22266 -21860 28186 -15940
rect 28585 -21860 34505 -15940
rect 34904 -21860 40824 -15940
rect 41223 -21860 47143 -15940
rect -47243 -28160 -41323 -22240
rect -40924 -28160 -35004 -22240
rect -34605 -28160 -28685 -22240
rect -28286 -28160 -22366 -22240
rect -21967 -28160 -16047 -22240
rect -15648 -28160 -9728 -22240
rect -9329 -28160 -3409 -22240
rect -3010 -28160 2910 -22240
rect 3309 -28160 9229 -22240
rect 9628 -28160 15548 -22240
rect 15947 -28160 21867 -22240
rect 22266 -28160 28186 -22240
rect 28585 -28160 34505 -22240
rect 34904 -28160 40824 -22240
rect 41223 -28160 47143 -22240
rect -47243 -34460 -41323 -28540
rect -40924 -34460 -35004 -28540
rect -34605 -34460 -28685 -28540
rect -28286 -34460 -22366 -28540
rect -21967 -34460 -16047 -28540
rect -15648 -34460 -9728 -28540
rect -9329 -34460 -3409 -28540
rect -3010 -34460 2910 -28540
rect 3309 -34460 9229 -28540
rect 9628 -34460 15548 -28540
rect 15947 -34460 21867 -28540
rect 22266 -34460 28186 -28540
rect 28585 -34460 34505 -28540
rect 34904 -34460 40824 -28540
rect 41223 -34460 47143 -28540
rect -47243 -40760 -41323 -34840
rect -40924 -40760 -35004 -34840
rect -34605 -40760 -28685 -34840
rect -28286 -40760 -22366 -34840
rect -21967 -40760 -16047 -34840
rect -15648 -40760 -9728 -34840
rect -9329 -40760 -3409 -34840
rect -3010 -40760 2910 -34840
rect 3309 -40760 9229 -34840
rect 9628 -40760 15548 -34840
rect 15947 -40760 21867 -34840
rect 22266 -40760 28186 -34840
rect 28585 -40760 34505 -34840
rect 34904 -40760 40824 -34840
rect 41223 -40760 47143 -34840
rect -47243 -47060 -41323 -41140
rect -40924 -47060 -35004 -41140
rect -34605 -47060 -28685 -41140
rect -28286 -47060 -22366 -41140
rect -21967 -47060 -16047 -41140
rect -15648 -47060 -9728 -41140
rect -9329 -47060 -3409 -41140
rect -3010 -47060 2910 -41140
rect 3309 -47060 9229 -41140
rect 9628 -47060 15548 -41140
rect 15947 -47060 21867 -41140
rect 22266 -47060 28186 -41140
rect 28585 -47060 34505 -41140
rect 34904 -47060 40824 -41140
rect 41223 -47060 47143 -41140
<< metal4 >>
rect -44335 47061 -44231 47250
rect -41215 47188 -41111 47250
rect -41215 47172 -41088 47188
rect -47244 47060 -41322 47061
rect -47244 41140 -47243 47060
rect -41323 41140 -41322 47060
rect -47244 41139 -41322 41140
rect -44335 40761 -44231 41139
rect -41215 41028 -41168 47172
rect -41104 41028 -41088 47172
rect -38016 47061 -37912 47250
rect -34896 47188 -34792 47250
rect -34896 47172 -34769 47188
rect -40925 47060 -35003 47061
rect -40925 41140 -40924 47060
rect -35004 41140 -35003 47060
rect -40925 41139 -35003 41140
rect -41215 41012 -41088 41028
rect -41215 40888 -41111 41012
rect -41215 40872 -41088 40888
rect -47244 40760 -41322 40761
rect -47244 34840 -47243 40760
rect -41323 34840 -41322 40760
rect -47244 34839 -41322 34840
rect -44335 34461 -44231 34839
rect -41215 34728 -41168 40872
rect -41104 34728 -41088 40872
rect -38016 40761 -37912 41139
rect -34896 41028 -34849 47172
rect -34785 41028 -34769 47172
rect -31697 47061 -31593 47250
rect -28577 47188 -28473 47250
rect -28577 47172 -28450 47188
rect -34606 47060 -28684 47061
rect -34606 41140 -34605 47060
rect -28685 41140 -28684 47060
rect -34606 41139 -28684 41140
rect -34896 41012 -34769 41028
rect -34896 40888 -34792 41012
rect -34896 40872 -34769 40888
rect -40925 40760 -35003 40761
rect -40925 34840 -40924 40760
rect -35004 34840 -35003 40760
rect -40925 34839 -35003 34840
rect -41215 34712 -41088 34728
rect -41215 34588 -41111 34712
rect -41215 34572 -41088 34588
rect -47244 34460 -41322 34461
rect -47244 28540 -47243 34460
rect -41323 28540 -41322 34460
rect -47244 28539 -41322 28540
rect -44335 28161 -44231 28539
rect -41215 28428 -41168 34572
rect -41104 28428 -41088 34572
rect -38016 34461 -37912 34839
rect -34896 34728 -34849 40872
rect -34785 34728 -34769 40872
rect -31697 40761 -31593 41139
rect -28577 41028 -28530 47172
rect -28466 41028 -28450 47172
rect -25378 47061 -25274 47250
rect -22258 47188 -22154 47250
rect -22258 47172 -22131 47188
rect -28287 47060 -22365 47061
rect -28287 41140 -28286 47060
rect -22366 41140 -22365 47060
rect -28287 41139 -22365 41140
rect -28577 41012 -28450 41028
rect -28577 40888 -28473 41012
rect -28577 40872 -28450 40888
rect -34606 40760 -28684 40761
rect -34606 34840 -34605 40760
rect -28685 34840 -28684 40760
rect -34606 34839 -28684 34840
rect -34896 34712 -34769 34728
rect -34896 34588 -34792 34712
rect -34896 34572 -34769 34588
rect -40925 34460 -35003 34461
rect -40925 28540 -40924 34460
rect -35004 28540 -35003 34460
rect -40925 28539 -35003 28540
rect -41215 28412 -41088 28428
rect -41215 28288 -41111 28412
rect -41215 28272 -41088 28288
rect -47244 28160 -41322 28161
rect -47244 22240 -47243 28160
rect -41323 22240 -41322 28160
rect -47244 22239 -41322 22240
rect -44335 21861 -44231 22239
rect -41215 22128 -41168 28272
rect -41104 22128 -41088 28272
rect -38016 28161 -37912 28539
rect -34896 28428 -34849 34572
rect -34785 28428 -34769 34572
rect -31697 34461 -31593 34839
rect -28577 34728 -28530 40872
rect -28466 34728 -28450 40872
rect -25378 40761 -25274 41139
rect -22258 41028 -22211 47172
rect -22147 41028 -22131 47172
rect -19059 47061 -18955 47250
rect -15939 47188 -15835 47250
rect -15939 47172 -15812 47188
rect -21968 47060 -16046 47061
rect -21968 41140 -21967 47060
rect -16047 41140 -16046 47060
rect -21968 41139 -16046 41140
rect -22258 41012 -22131 41028
rect -22258 40888 -22154 41012
rect -22258 40872 -22131 40888
rect -28287 40760 -22365 40761
rect -28287 34840 -28286 40760
rect -22366 34840 -22365 40760
rect -28287 34839 -22365 34840
rect -28577 34712 -28450 34728
rect -28577 34588 -28473 34712
rect -28577 34572 -28450 34588
rect -34606 34460 -28684 34461
rect -34606 28540 -34605 34460
rect -28685 28540 -28684 34460
rect -34606 28539 -28684 28540
rect -34896 28412 -34769 28428
rect -34896 28288 -34792 28412
rect -34896 28272 -34769 28288
rect -40925 28160 -35003 28161
rect -40925 22240 -40924 28160
rect -35004 22240 -35003 28160
rect -40925 22239 -35003 22240
rect -41215 22112 -41088 22128
rect -41215 21988 -41111 22112
rect -41215 21972 -41088 21988
rect -47244 21860 -41322 21861
rect -47244 15940 -47243 21860
rect -41323 15940 -41322 21860
rect -47244 15939 -41322 15940
rect -44335 15561 -44231 15939
rect -41215 15828 -41168 21972
rect -41104 15828 -41088 21972
rect -38016 21861 -37912 22239
rect -34896 22128 -34849 28272
rect -34785 22128 -34769 28272
rect -31697 28161 -31593 28539
rect -28577 28428 -28530 34572
rect -28466 28428 -28450 34572
rect -25378 34461 -25274 34839
rect -22258 34728 -22211 40872
rect -22147 34728 -22131 40872
rect -19059 40761 -18955 41139
rect -15939 41028 -15892 47172
rect -15828 41028 -15812 47172
rect -12740 47061 -12636 47250
rect -9620 47188 -9516 47250
rect -9620 47172 -9493 47188
rect -15649 47060 -9727 47061
rect -15649 41140 -15648 47060
rect -9728 41140 -9727 47060
rect -15649 41139 -9727 41140
rect -15939 41012 -15812 41028
rect -15939 40888 -15835 41012
rect -15939 40872 -15812 40888
rect -21968 40760 -16046 40761
rect -21968 34840 -21967 40760
rect -16047 34840 -16046 40760
rect -21968 34839 -16046 34840
rect -22258 34712 -22131 34728
rect -22258 34588 -22154 34712
rect -22258 34572 -22131 34588
rect -28287 34460 -22365 34461
rect -28287 28540 -28286 34460
rect -22366 28540 -22365 34460
rect -28287 28539 -22365 28540
rect -28577 28412 -28450 28428
rect -28577 28288 -28473 28412
rect -28577 28272 -28450 28288
rect -34606 28160 -28684 28161
rect -34606 22240 -34605 28160
rect -28685 22240 -28684 28160
rect -34606 22239 -28684 22240
rect -34896 22112 -34769 22128
rect -34896 21988 -34792 22112
rect -34896 21972 -34769 21988
rect -40925 21860 -35003 21861
rect -40925 15940 -40924 21860
rect -35004 15940 -35003 21860
rect -40925 15939 -35003 15940
rect -41215 15812 -41088 15828
rect -41215 15688 -41111 15812
rect -41215 15672 -41088 15688
rect -47244 15560 -41322 15561
rect -47244 9640 -47243 15560
rect -41323 9640 -41322 15560
rect -47244 9639 -41322 9640
rect -44335 9261 -44231 9639
rect -41215 9528 -41168 15672
rect -41104 9528 -41088 15672
rect -38016 15561 -37912 15939
rect -34896 15828 -34849 21972
rect -34785 15828 -34769 21972
rect -31697 21861 -31593 22239
rect -28577 22128 -28530 28272
rect -28466 22128 -28450 28272
rect -25378 28161 -25274 28539
rect -22258 28428 -22211 34572
rect -22147 28428 -22131 34572
rect -19059 34461 -18955 34839
rect -15939 34728 -15892 40872
rect -15828 34728 -15812 40872
rect -12740 40761 -12636 41139
rect -9620 41028 -9573 47172
rect -9509 41028 -9493 47172
rect -6421 47061 -6317 47250
rect -3301 47188 -3197 47250
rect -3301 47172 -3174 47188
rect -9330 47060 -3408 47061
rect -9330 41140 -9329 47060
rect -3409 41140 -3408 47060
rect -9330 41139 -3408 41140
rect -9620 41012 -9493 41028
rect -9620 40888 -9516 41012
rect -9620 40872 -9493 40888
rect -15649 40760 -9727 40761
rect -15649 34840 -15648 40760
rect -9728 34840 -9727 40760
rect -15649 34839 -9727 34840
rect -15939 34712 -15812 34728
rect -15939 34588 -15835 34712
rect -15939 34572 -15812 34588
rect -21968 34460 -16046 34461
rect -21968 28540 -21967 34460
rect -16047 28540 -16046 34460
rect -21968 28539 -16046 28540
rect -22258 28412 -22131 28428
rect -22258 28288 -22154 28412
rect -22258 28272 -22131 28288
rect -28287 28160 -22365 28161
rect -28287 22240 -28286 28160
rect -22366 22240 -22365 28160
rect -28287 22239 -22365 22240
rect -28577 22112 -28450 22128
rect -28577 21988 -28473 22112
rect -28577 21972 -28450 21988
rect -34606 21860 -28684 21861
rect -34606 15940 -34605 21860
rect -28685 15940 -28684 21860
rect -34606 15939 -28684 15940
rect -34896 15812 -34769 15828
rect -34896 15688 -34792 15812
rect -34896 15672 -34769 15688
rect -40925 15560 -35003 15561
rect -40925 9640 -40924 15560
rect -35004 9640 -35003 15560
rect -40925 9639 -35003 9640
rect -41215 9512 -41088 9528
rect -41215 9388 -41111 9512
rect -41215 9372 -41088 9388
rect -47244 9260 -41322 9261
rect -47244 3340 -47243 9260
rect -41323 3340 -41322 9260
rect -47244 3339 -41322 3340
rect -44335 2961 -44231 3339
rect -41215 3228 -41168 9372
rect -41104 3228 -41088 9372
rect -38016 9261 -37912 9639
rect -34896 9528 -34849 15672
rect -34785 9528 -34769 15672
rect -31697 15561 -31593 15939
rect -28577 15828 -28530 21972
rect -28466 15828 -28450 21972
rect -25378 21861 -25274 22239
rect -22258 22128 -22211 28272
rect -22147 22128 -22131 28272
rect -19059 28161 -18955 28539
rect -15939 28428 -15892 34572
rect -15828 28428 -15812 34572
rect -12740 34461 -12636 34839
rect -9620 34728 -9573 40872
rect -9509 34728 -9493 40872
rect -6421 40761 -6317 41139
rect -3301 41028 -3254 47172
rect -3190 41028 -3174 47172
rect -102 47061 2 47250
rect 3018 47188 3122 47250
rect 3018 47172 3145 47188
rect -3011 47060 2911 47061
rect -3011 41140 -3010 47060
rect 2910 41140 2911 47060
rect -3011 41139 2911 41140
rect -3301 41012 -3174 41028
rect -3301 40888 -3197 41012
rect -3301 40872 -3174 40888
rect -9330 40760 -3408 40761
rect -9330 34840 -9329 40760
rect -3409 34840 -3408 40760
rect -9330 34839 -3408 34840
rect -9620 34712 -9493 34728
rect -9620 34588 -9516 34712
rect -9620 34572 -9493 34588
rect -15649 34460 -9727 34461
rect -15649 28540 -15648 34460
rect -9728 28540 -9727 34460
rect -15649 28539 -9727 28540
rect -15939 28412 -15812 28428
rect -15939 28288 -15835 28412
rect -15939 28272 -15812 28288
rect -21968 28160 -16046 28161
rect -21968 22240 -21967 28160
rect -16047 22240 -16046 28160
rect -21968 22239 -16046 22240
rect -22258 22112 -22131 22128
rect -22258 21988 -22154 22112
rect -22258 21972 -22131 21988
rect -28287 21860 -22365 21861
rect -28287 15940 -28286 21860
rect -22366 15940 -22365 21860
rect -28287 15939 -22365 15940
rect -28577 15812 -28450 15828
rect -28577 15688 -28473 15812
rect -28577 15672 -28450 15688
rect -34606 15560 -28684 15561
rect -34606 9640 -34605 15560
rect -28685 9640 -28684 15560
rect -34606 9639 -28684 9640
rect -34896 9512 -34769 9528
rect -34896 9388 -34792 9512
rect -34896 9372 -34769 9388
rect -40925 9260 -35003 9261
rect -40925 3340 -40924 9260
rect -35004 3340 -35003 9260
rect -40925 3339 -35003 3340
rect -41215 3212 -41088 3228
rect -41215 3088 -41111 3212
rect -41215 3072 -41088 3088
rect -47244 2960 -41322 2961
rect -47244 -2960 -47243 2960
rect -41323 -2960 -41322 2960
rect -47244 -2961 -41322 -2960
rect -44335 -3339 -44231 -2961
rect -41215 -3072 -41168 3072
rect -41104 -3072 -41088 3072
rect -38016 2961 -37912 3339
rect -34896 3228 -34849 9372
rect -34785 3228 -34769 9372
rect -31697 9261 -31593 9639
rect -28577 9528 -28530 15672
rect -28466 9528 -28450 15672
rect -25378 15561 -25274 15939
rect -22258 15828 -22211 21972
rect -22147 15828 -22131 21972
rect -19059 21861 -18955 22239
rect -15939 22128 -15892 28272
rect -15828 22128 -15812 28272
rect -12740 28161 -12636 28539
rect -9620 28428 -9573 34572
rect -9509 28428 -9493 34572
rect -6421 34461 -6317 34839
rect -3301 34728 -3254 40872
rect -3190 34728 -3174 40872
rect -102 40761 2 41139
rect 3018 41028 3065 47172
rect 3129 41028 3145 47172
rect 6217 47061 6321 47250
rect 9337 47188 9441 47250
rect 9337 47172 9464 47188
rect 3308 47060 9230 47061
rect 3308 41140 3309 47060
rect 9229 41140 9230 47060
rect 3308 41139 9230 41140
rect 3018 41012 3145 41028
rect 3018 40888 3122 41012
rect 3018 40872 3145 40888
rect -3011 40760 2911 40761
rect -3011 34840 -3010 40760
rect 2910 34840 2911 40760
rect -3011 34839 2911 34840
rect -3301 34712 -3174 34728
rect -3301 34588 -3197 34712
rect -3301 34572 -3174 34588
rect -9330 34460 -3408 34461
rect -9330 28540 -9329 34460
rect -3409 28540 -3408 34460
rect -9330 28539 -3408 28540
rect -9620 28412 -9493 28428
rect -9620 28288 -9516 28412
rect -9620 28272 -9493 28288
rect -15649 28160 -9727 28161
rect -15649 22240 -15648 28160
rect -9728 22240 -9727 28160
rect -15649 22239 -9727 22240
rect -15939 22112 -15812 22128
rect -15939 21988 -15835 22112
rect -15939 21972 -15812 21988
rect -21968 21860 -16046 21861
rect -21968 15940 -21967 21860
rect -16047 15940 -16046 21860
rect -21968 15939 -16046 15940
rect -22258 15812 -22131 15828
rect -22258 15688 -22154 15812
rect -22258 15672 -22131 15688
rect -28287 15560 -22365 15561
rect -28287 9640 -28286 15560
rect -22366 9640 -22365 15560
rect -28287 9639 -22365 9640
rect -28577 9512 -28450 9528
rect -28577 9388 -28473 9512
rect -28577 9372 -28450 9388
rect -34606 9260 -28684 9261
rect -34606 3340 -34605 9260
rect -28685 3340 -28684 9260
rect -34606 3339 -28684 3340
rect -34896 3212 -34769 3228
rect -34896 3088 -34792 3212
rect -34896 3072 -34769 3088
rect -40925 2960 -35003 2961
rect -40925 -2960 -40924 2960
rect -35004 -2960 -35003 2960
rect -40925 -2961 -35003 -2960
rect -41215 -3088 -41088 -3072
rect -41215 -3212 -41111 -3088
rect -41215 -3228 -41088 -3212
rect -47244 -3340 -41322 -3339
rect -47244 -9260 -47243 -3340
rect -41323 -9260 -41322 -3340
rect -47244 -9261 -41322 -9260
rect -44335 -9639 -44231 -9261
rect -41215 -9372 -41168 -3228
rect -41104 -9372 -41088 -3228
rect -38016 -3339 -37912 -2961
rect -34896 -3072 -34849 3072
rect -34785 -3072 -34769 3072
rect -31697 2961 -31593 3339
rect -28577 3228 -28530 9372
rect -28466 3228 -28450 9372
rect -25378 9261 -25274 9639
rect -22258 9528 -22211 15672
rect -22147 9528 -22131 15672
rect -19059 15561 -18955 15939
rect -15939 15828 -15892 21972
rect -15828 15828 -15812 21972
rect -12740 21861 -12636 22239
rect -9620 22128 -9573 28272
rect -9509 22128 -9493 28272
rect -6421 28161 -6317 28539
rect -3301 28428 -3254 34572
rect -3190 28428 -3174 34572
rect -102 34461 2 34839
rect 3018 34728 3065 40872
rect 3129 34728 3145 40872
rect 6217 40761 6321 41139
rect 9337 41028 9384 47172
rect 9448 41028 9464 47172
rect 12536 47061 12640 47250
rect 15656 47188 15760 47250
rect 15656 47172 15783 47188
rect 9627 47060 15549 47061
rect 9627 41140 9628 47060
rect 15548 41140 15549 47060
rect 9627 41139 15549 41140
rect 9337 41012 9464 41028
rect 9337 40888 9441 41012
rect 9337 40872 9464 40888
rect 3308 40760 9230 40761
rect 3308 34840 3309 40760
rect 9229 34840 9230 40760
rect 3308 34839 9230 34840
rect 3018 34712 3145 34728
rect 3018 34588 3122 34712
rect 3018 34572 3145 34588
rect -3011 34460 2911 34461
rect -3011 28540 -3010 34460
rect 2910 28540 2911 34460
rect -3011 28539 2911 28540
rect -3301 28412 -3174 28428
rect -3301 28288 -3197 28412
rect -3301 28272 -3174 28288
rect -9330 28160 -3408 28161
rect -9330 22240 -9329 28160
rect -3409 22240 -3408 28160
rect -9330 22239 -3408 22240
rect -9620 22112 -9493 22128
rect -9620 21988 -9516 22112
rect -9620 21972 -9493 21988
rect -15649 21860 -9727 21861
rect -15649 15940 -15648 21860
rect -9728 15940 -9727 21860
rect -15649 15939 -9727 15940
rect -15939 15812 -15812 15828
rect -15939 15688 -15835 15812
rect -15939 15672 -15812 15688
rect -21968 15560 -16046 15561
rect -21968 9640 -21967 15560
rect -16047 9640 -16046 15560
rect -21968 9639 -16046 9640
rect -22258 9512 -22131 9528
rect -22258 9388 -22154 9512
rect -22258 9372 -22131 9388
rect -28287 9260 -22365 9261
rect -28287 3340 -28286 9260
rect -22366 3340 -22365 9260
rect -28287 3339 -22365 3340
rect -28577 3212 -28450 3228
rect -28577 3088 -28473 3212
rect -28577 3072 -28450 3088
rect -34606 2960 -28684 2961
rect -34606 -2960 -34605 2960
rect -28685 -2960 -28684 2960
rect -34606 -2961 -28684 -2960
rect -34896 -3088 -34769 -3072
rect -34896 -3212 -34792 -3088
rect -34896 -3228 -34769 -3212
rect -40925 -3340 -35003 -3339
rect -40925 -9260 -40924 -3340
rect -35004 -9260 -35003 -3340
rect -40925 -9261 -35003 -9260
rect -41215 -9388 -41088 -9372
rect -41215 -9512 -41111 -9388
rect -41215 -9528 -41088 -9512
rect -47244 -9640 -41322 -9639
rect -47244 -15560 -47243 -9640
rect -41323 -15560 -41322 -9640
rect -47244 -15561 -41322 -15560
rect -44335 -15939 -44231 -15561
rect -41215 -15672 -41168 -9528
rect -41104 -15672 -41088 -9528
rect -38016 -9639 -37912 -9261
rect -34896 -9372 -34849 -3228
rect -34785 -9372 -34769 -3228
rect -31697 -3339 -31593 -2961
rect -28577 -3072 -28530 3072
rect -28466 -3072 -28450 3072
rect -25378 2961 -25274 3339
rect -22258 3228 -22211 9372
rect -22147 3228 -22131 9372
rect -19059 9261 -18955 9639
rect -15939 9528 -15892 15672
rect -15828 9528 -15812 15672
rect -12740 15561 -12636 15939
rect -9620 15828 -9573 21972
rect -9509 15828 -9493 21972
rect -6421 21861 -6317 22239
rect -3301 22128 -3254 28272
rect -3190 22128 -3174 28272
rect -102 28161 2 28539
rect 3018 28428 3065 34572
rect 3129 28428 3145 34572
rect 6217 34461 6321 34839
rect 9337 34728 9384 40872
rect 9448 34728 9464 40872
rect 12536 40761 12640 41139
rect 15656 41028 15703 47172
rect 15767 41028 15783 47172
rect 18855 47061 18959 47250
rect 21975 47188 22079 47250
rect 21975 47172 22102 47188
rect 15946 47060 21868 47061
rect 15946 41140 15947 47060
rect 21867 41140 21868 47060
rect 15946 41139 21868 41140
rect 15656 41012 15783 41028
rect 15656 40888 15760 41012
rect 15656 40872 15783 40888
rect 9627 40760 15549 40761
rect 9627 34840 9628 40760
rect 15548 34840 15549 40760
rect 9627 34839 15549 34840
rect 9337 34712 9464 34728
rect 9337 34588 9441 34712
rect 9337 34572 9464 34588
rect 3308 34460 9230 34461
rect 3308 28540 3309 34460
rect 9229 28540 9230 34460
rect 3308 28539 9230 28540
rect 3018 28412 3145 28428
rect 3018 28288 3122 28412
rect 3018 28272 3145 28288
rect -3011 28160 2911 28161
rect -3011 22240 -3010 28160
rect 2910 22240 2911 28160
rect -3011 22239 2911 22240
rect -3301 22112 -3174 22128
rect -3301 21988 -3197 22112
rect -3301 21972 -3174 21988
rect -9330 21860 -3408 21861
rect -9330 15940 -9329 21860
rect -3409 15940 -3408 21860
rect -9330 15939 -3408 15940
rect -9620 15812 -9493 15828
rect -9620 15688 -9516 15812
rect -9620 15672 -9493 15688
rect -15649 15560 -9727 15561
rect -15649 9640 -15648 15560
rect -9728 9640 -9727 15560
rect -15649 9639 -9727 9640
rect -15939 9512 -15812 9528
rect -15939 9388 -15835 9512
rect -15939 9372 -15812 9388
rect -21968 9260 -16046 9261
rect -21968 3340 -21967 9260
rect -16047 3340 -16046 9260
rect -21968 3339 -16046 3340
rect -22258 3212 -22131 3228
rect -22258 3088 -22154 3212
rect -22258 3072 -22131 3088
rect -28287 2960 -22365 2961
rect -28287 -2960 -28286 2960
rect -22366 -2960 -22365 2960
rect -28287 -2961 -22365 -2960
rect -28577 -3088 -28450 -3072
rect -28577 -3212 -28473 -3088
rect -28577 -3228 -28450 -3212
rect -34606 -3340 -28684 -3339
rect -34606 -9260 -34605 -3340
rect -28685 -9260 -28684 -3340
rect -34606 -9261 -28684 -9260
rect -34896 -9388 -34769 -9372
rect -34896 -9512 -34792 -9388
rect -34896 -9528 -34769 -9512
rect -40925 -9640 -35003 -9639
rect -40925 -15560 -40924 -9640
rect -35004 -15560 -35003 -9640
rect -40925 -15561 -35003 -15560
rect -41215 -15688 -41088 -15672
rect -41215 -15812 -41111 -15688
rect -41215 -15828 -41088 -15812
rect -47244 -15940 -41322 -15939
rect -47244 -21860 -47243 -15940
rect -41323 -21860 -41322 -15940
rect -47244 -21861 -41322 -21860
rect -44335 -22239 -44231 -21861
rect -41215 -21972 -41168 -15828
rect -41104 -21972 -41088 -15828
rect -38016 -15939 -37912 -15561
rect -34896 -15672 -34849 -9528
rect -34785 -15672 -34769 -9528
rect -31697 -9639 -31593 -9261
rect -28577 -9372 -28530 -3228
rect -28466 -9372 -28450 -3228
rect -25378 -3339 -25274 -2961
rect -22258 -3072 -22211 3072
rect -22147 -3072 -22131 3072
rect -19059 2961 -18955 3339
rect -15939 3228 -15892 9372
rect -15828 3228 -15812 9372
rect -12740 9261 -12636 9639
rect -9620 9528 -9573 15672
rect -9509 9528 -9493 15672
rect -6421 15561 -6317 15939
rect -3301 15828 -3254 21972
rect -3190 15828 -3174 21972
rect -102 21861 2 22239
rect 3018 22128 3065 28272
rect 3129 22128 3145 28272
rect 6217 28161 6321 28539
rect 9337 28428 9384 34572
rect 9448 28428 9464 34572
rect 12536 34461 12640 34839
rect 15656 34728 15703 40872
rect 15767 34728 15783 40872
rect 18855 40761 18959 41139
rect 21975 41028 22022 47172
rect 22086 41028 22102 47172
rect 25174 47061 25278 47250
rect 28294 47188 28398 47250
rect 28294 47172 28421 47188
rect 22265 47060 28187 47061
rect 22265 41140 22266 47060
rect 28186 41140 28187 47060
rect 22265 41139 28187 41140
rect 21975 41012 22102 41028
rect 21975 40888 22079 41012
rect 21975 40872 22102 40888
rect 15946 40760 21868 40761
rect 15946 34840 15947 40760
rect 21867 34840 21868 40760
rect 15946 34839 21868 34840
rect 15656 34712 15783 34728
rect 15656 34588 15760 34712
rect 15656 34572 15783 34588
rect 9627 34460 15549 34461
rect 9627 28540 9628 34460
rect 15548 28540 15549 34460
rect 9627 28539 15549 28540
rect 9337 28412 9464 28428
rect 9337 28288 9441 28412
rect 9337 28272 9464 28288
rect 3308 28160 9230 28161
rect 3308 22240 3309 28160
rect 9229 22240 9230 28160
rect 3308 22239 9230 22240
rect 3018 22112 3145 22128
rect 3018 21988 3122 22112
rect 3018 21972 3145 21988
rect -3011 21860 2911 21861
rect -3011 15940 -3010 21860
rect 2910 15940 2911 21860
rect -3011 15939 2911 15940
rect -3301 15812 -3174 15828
rect -3301 15688 -3197 15812
rect -3301 15672 -3174 15688
rect -9330 15560 -3408 15561
rect -9330 9640 -9329 15560
rect -3409 9640 -3408 15560
rect -9330 9639 -3408 9640
rect -9620 9512 -9493 9528
rect -9620 9388 -9516 9512
rect -9620 9372 -9493 9388
rect -15649 9260 -9727 9261
rect -15649 3340 -15648 9260
rect -9728 3340 -9727 9260
rect -15649 3339 -9727 3340
rect -15939 3212 -15812 3228
rect -15939 3088 -15835 3212
rect -15939 3072 -15812 3088
rect -21968 2960 -16046 2961
rect -21968 -2960 -21967 2960
rect -16047 -2960 -16046 2960
rect -21968 -2961 -16046 -2960
rect -22258 -3088 -22131 -3072
rect -22258 -3212 -22154 -3088
rect -22258 -3228 -22131 -3212
rect -28287 -3340 -22365 -3339
rect -28287 -9260 -28286 -3340
rect -22366 -9260 -22365 -3340
rect -28287 -9261 -22365 -9260
rect -28577 -9388 -28450 -9372
rect -28577 -9512 -28473 -9388
rect -28577 -9528 -28450 -9512
rect -34606 -9640 -28684 -9639
rect -34606 -15560 -34605 -9640
rect -28685 -15560 -28684 -9640
rect -34606 -15561 -28684 -15560
rect -34896 -15688 -34769 -15672
rect -34896 -15812 -34792 -15688
rect -34896 -15828 -34769 -15812
rect -40925 -15940 -35003 -15939
rect -40925 -21860 -40924 -15940
rect -35004 -21860 -35003 -15940
rect -40925 -21861 -35003 -21860
rect -41215 -21988 -41088 -21972
rect -41215 -22112 -41111 -21988
rect -41215 -22128 -41088 -22112
rect -47244 -22240 -41322 -22239
rect -47244 -28160 -47243 -22240
rect -41323 -28160 -41322 -22240
rect -47244 -28161 -41322 -28160
rect -44335 -28539 -44231 -28161
rect -41215 -28272 -41168 -22128
rect -41104 -28272 -41088 -22128
rect -38016 -22239 -37912 -21861
rect -34896 -21972 -34849 -15828
rect -34785 -21972 -34769 -15828
rect -31697 -15939 -31593 -15561
rect -28577 -15672 -28530 -9528
rect -28466 -15672 -28450 -9528
rect -25378 -9639 -25274 -9261
rect -22258 -9372 -22211 -3228
rect -22147 -9372 -22131 -3228
rect -19059 -3339 -18955 -2961
rect -15939 -3072 -15892 3072
rect -15828 -3072 -15812 3072
rect -12740 2961 -12636 3339
rect -9620 3228 -9573 9372
rect -9509 3228 -9493 9372
rect -6421 9261 -6317 9639
rect -3301 9528 -3254 15672
rect -3190 9528 -3174 15672
rect -102 15561 2 15939
rect 3018 15828 3065 21972
rect 3129 15828 3145 21972
rect 6217 21861 6321 22239
rect 9337 22128 9384 28272
rect 9448 22128 9464 28272
rect 12536 28161 12640 28539
rect 15656 28428 15703 34572
rect 15767 28428 15783 34572
rect 18855 34461 18959 34839
rect 21975 34728 22022 40872
rect 22086 34728 22102 40872
rect 25174 40761 25278 41139
rect 28294 41028 28341 47172
rect 28405 41028 28421 47172
rect 31493 47061 31597 47250
rect 34613 47188 34717 47250
rect 34613 47172 34740 47188
rect 28584 47060 34506 47061
rect 28584 41140 28585 47060
rect 34505 41140 34506 47060
rect 28584 41139 34506 41140
rect 28294 41012 28421 41028
rect 28294 40888 28398 41012
rect 28294 40872 28421 40888
rect 22265 40760 28187 40761
rect 22265 34840 22266 40760
rect 28186 34840 28187 40760
rect 22265 34839 28187 34840
rect 21975 34712 22102 34728
rect 21975 34588 22079 34712
rect 21975 34572 22102 34588
rect 15946 34460 21868 34461
rect 15946 28540 15947 34460
rect 21867 28540 21868 34460
rect 15946 28539 21868 28540
rect 15656 28412 15783 28428
rect 15656 28288 15760 28412
rect 15656 28272 15783 28288
rect 9627 28160 15549 28161
rect 9627 22240 9628 28160
rect 15548 22240 15549 28160
rect 9627 22239 15549 22240
rect 9337 22112 9464 22128
rect 9337 21988 9441 22112
rect 9337 21972 9464 21988
rect 3308 21860 9230 21861
rect 3308 15940 3309 21860
rect 9229 15940 9230 21860
rect 3308 15939 9230 15940
rect 3018 15812 3145 15828
rect 3018 15688 3122 15812
rect 3018 15672 3145 15688
rect -3011 15560 2911 15561
rect -3011 9640 -3010 15560
rect 2910 9640 2911 15560
rect -3011 9639 2911 9640
rect -3301 9512 -3174 9528
rect -3301 9388 -3197 9512
rect -3301 9372 -3174 9388
rect -9330 9260 -3408 9261
rect -9330 3340 -9329 9260
rect -3409 3340 -3408 9260
rect -9330 3339 -3408 3340
rect -9620 3212 -9493 3228
rect -9620 3088 -9516 3212
rect -9620 3072 -9493 3088
rect -15649 2960 -9727 2961
rect -15649 -2960 -15648 2960
rect -9728 -2960 -9727 2960
rect -15649 -2961 -9727 -2960
rect -15939 -3088 -15812 -3072
rect -15939 -3212 -15835 -3088
rect -15939 -3228 -15812 -3212
rect -21968 -3340 -16046 -3339
rect -21968 -9260 -21967 -3340
rect -16047 -9260 -16046 -3340
rect -21968 -9261 -16046 -9260
rect -22258 -9388 -22131 -9372
rect -22258 -9512 -22154 -9388
rect -22258 -9528 -22131 -9512
rect -28287 -9640 -22365 -9639
rect -28287 -15560 -28286 -9640
rect -22366 -15560 -22365 -9640
rect -28287 -15561 -22365 -15560
rect -28577 -15688 -28450 -15672
rect -28577 -15812 -28473 -15688
rect -28577 -15828 -28450 -15812
rect -34606 -15940 -28684 -15939
rect -34606 -21860 -34605 -15940
rect -28685 -21860 -28684 -15940
rect -34606 -21861 -28684 -21860
rect -34896 -21988 -34769 -21972
rect -34896 -22112 -34792 -21988
rect -34896 -22128 -34769 -22112
rect -40925 -22240 -35003 -22239
rect -40925 -28160 -40924 -22240
rect -35004 -28160 -35003 -22240
rect -40925 -28161 -35003 -28160
rect -41215 -28288 -41088 -28272
rect -41215 -28412 -41111 -28288
rect -41215 -28428 -41088 -28412
rect -47244 -28540 -41322 -28539
rect -47244 -34460 -47243 -28540
rect -41323 -34460 -41322 -28540
rect -47244 -34461 -41322 -34460
rect -44335 -34839 -44231 -34461
rect -41215 -34572 -41168 -28428
rect -41104 -34572 -41088 -28428
rect -38016 -28539 -37912 -28161
rect -34896 -28272 -34849 -22128
rect -34785 -28272 -34769 -22128
rect -31697 -22239 -31593 -21861
rect -28577 -21972 -28530 -15828
rect -28466 -21972 -28450 -15828
rect -25378 -15939 -25274 -15561
rect -22258 -15672 -22211 -9528
rect -22147 -15672 -22131 -9528
rect -19059 -9639 -18955 -9261
rect -15939 -9372 -15892 -3228
rect -15828 -9372 -15812 -3228
rect -12740 -3339 -12636 -2961
rect -9620 -3072 -9573 3072
rect -9509 -3072 -9493 3072
rect -6421 2961 -6317 3339
rect -3301 3228 -3254 9372
rect -3190 3228 -3174 9372
rect -102 9261 2 9639
rect 3018 9528 3065 15672
rect 3129 9528 3145 15672
rect 6217 15561 6321 15939
rect 9337 15828 9384 21972
rect 9448 15828 9464 21972
rect 12536 21861 12640 22239
rect 15656 22128 15703 28272
rect 15767 22128 15783 28272
rect 18855 28161 18959 28539
rect 21975 28428 22022 34572
rect 22086 28428 22102 34572
rect 25174 34461 25278 34839
rect 28294 34728 28341 40872
rect 28405 34728 28421 40872
rect 31493 40761 31597 41139
rect 34613 41028 34660 47172
rect 34724 41028 34740 47172
rect 37812 47061 37916 47250
rect 40932 47188 41036 47250
rect 40932 47172 41059 47188
rect 34903 47060 40825 47061
rect 34903 41140 34904 47060
rect 40824 41140 40825 47060
rect 34903 41139 40825 41140
rect 34613 41012 34740 41028
rect 34613 40888 34717 41012
rect 34613 40872 34740 40888
rect 28584 40760 34506 40761
rect 28584 34840 28585 40760
rect 34505 34840 34506 40760
rect 28584 34839 34506 34840
rect 28294 34712 28421 34728
rect 28294 34588 28398 34712
rect 28294 34572 28421 34588
rect 22265 34460 28187 34461
rect 22265 28540 22266 34460
rect 28186 28540 28187 34460
rect 22265 28539 28187 28540
rect 21975 28412 22102 28428
rect 21975 28288 22079 28412
rect 21975 28272 22102 28288
rect 15946 28160 21868 28161
rect 15946 22240 15947 28160
rect 21867 22240 21868 28160
rect 15946 22239 21868 22240
rect 15656 22112 15783 22128
rect 15656 21988 15760 22112
rect 15656 21972 15783 21988
rect 9627 21860 15549 21861
rect 9627 15940 9628 21860
rect 15548 15940 15549 21860
rect 9627 15939 15549 15940
rect 9337 15812 9464 15828
rect 9337 15688 9441 15812
rect 9337 15672 9464 15688
rect 3308 15560 9230 15561
rect 3308 9640 3309 15560
rect 9229 9640 9230 15560
rect 3308 9639 9230 9640
rect 3018 9512 3145 9528
rect 3018 9388 3122 9512
rect 3018 9372 3145 9388
rect -3011 9260 2911 9261
rect -3011 3340 -3010 9260
rect 2910 3340 2911 9260
rect -3011 3339 2911 3340
rect -3301 3212 -3174 3228
rect -3301 3088 -3197 3212
rect -3301 3072 -3174 3088
rect -9330 2960 -3408 2961
rect -9330 -2960 -9329 2960
rect -3409 -2960 -3408 2960
rect -9330 -2961 -3408 -2960
rect -9620 -3088 -9493 -3072
rect -9620 -3212 -9516 -3088
rect -9620 -3228 -9493 -3212
rect -15649 -3340 -9727 -3339
rect -15649 -9260 -15648 -3340
rect -9728 -9260 -9727 -3340
rect -15649 -9261 -9727 -9260
rect -15939 -9388 -15812 -9372
rect -15939 -9512 -15835 -9388
rect -15939 -9528 -15812 -9512
rect -21968 -9640 -16046 -9639
rect -21968 -15560 -21967 -9640
rect -16047 -15560 -16046 -9640
rect -21968 -15561 -16046 -15560
rect -22258 -15688 -22131 -15672
rect -22258 -15812 -22154 -15688
rect -22258 -15828 -22131 -15812
rect -28287 -15940 -22365 -15939
rect -28287 -21860 -28286 -15940
rect -22366 -21860 -22365 -15940
rect -28287 -21861 -22365 -21860
rect -28577 -21988 -28450 -21972
rect -28577 -22112 -28473 -21988
rect -28577 -22128 -28450 -22112
rect -34606 -22240 -28684 -22239
rect -34606 -28160 -34605 -22240
rect -28685 -28160 -28684 -22240
rect -34606 -28161 -28684 -28160
rect -34896 -28288 -34769 -28272
rect -34896 -28412 -34792 -28288
rect -34896 -28428 -34769 -28412
rect -40925 -28540 -35003 -28539
rect -40925 -34460 -40924 -28540
rect -35004 -34460 -35003 -28540
rect -40925 -34461 -35003 -34460
rect -41215 -34588 -41088 -34572
rect -41215 -34712 -41111 -34588
rect -41215 -34728 -41088 -34712
rect -47244 -34840 -41322 -34839
rect -47244 -40760 -47243 -34840
rect -41323 -40760 -41322 -34840
rect -47244 -40761 -41322 -40760
rect -44335 -41139 -44231 -40761
rect -41215 -40872 -41168 -34728
rect -41104 -40872 -41088 -34728
rect -38016 -34839 -37912 -34461
rect -34896 -34572 -34849 -28428
rect -34785 -34572 -34769 -28428
rect -31697 -28539 -31593 -28161
rect -28577 -28272 -28530 -22128
rect -28466 -28272 -28450 -22128
rect -25378 -22239 -25274 -21861
rect -22258 -21972 -22211 -15828
rect -22147 -21972 -22131 -15828
rect -19059 -15939 -18955 -15561
rect -15939 -15672 -15892 -9528
rect -15828 -15672 -15812 -9528
rect -12740 -9639 -12636 -9261
rect -9620 -9372 -9573 -3228
rect -9509 -9372 -9493 -3228
rect -6421 -3339 -6317 -2961
rect -3301 -3072 -3254 3072
rect -3190 -3072 -3174 3072
rect -102 2961 2 3339
rect 3018 3228 3065 9372
rect 3129 3228 3145 9372
rect 6217 9261 6321 9639
rect 9337 9528 9384 15672
rect 9448 9528 9464 15672
rect 12536 15561 12640 15939
rect 15656 15828 15703 21972
rect 15767 15828 15783 21972
rect 18855 21861 18959 22239
rect 21975 22128 22022 28272
rect 22086 22128 22102 28272
rect 25174 28161 25278 28539
rect 28294 28428 28341 34572
rect 28405 28428 28421 34572
rect 31493 34461 31597 34839
rect 34613 34728 34660 40872
rect 34724 34728 34740 40872
rect 37812 40761 37916 41139
rect 40932 41028 40979 47172
rect 41043 41028 41059 47172
rect 44131 47061 44235 47250
rect 47251 47188 47355 47250
rect 47251 47172 47378 47188
rect 41222 47060 47144 47061
rect 41222 41140 41223 47060
rect 47143 41140 47144 47060
rect 41222 41139 47144 41140
rect 40932 41012 41059 41028
rect 40932 40888 41036 41012
rect 40932 40872 41059 40888
rect 34903 40760 40825 40761
rect 34903 34840 34904 40760
rect 40824 34840 40825 40760
rect 34903 34839 40825 34840
rect 34613 34712 34740 34728
rect 34613 34588 34717 34712
rect 34613 34572 34740 34588
rect 28584 34460 34506 34461
rect 28584 28540 28585 34460
rect 34505 28540 34506 34460
rect 28584 28539 34506 28540
rect 28294 28412 28421 28428
rect 28294 28288 28398 28412
rect 28294 28272 28421 28288
rect 22265 28160 28187 28161
rect 22265 22240 22266 28160
rect 28186 22240 28187 28160
rect 22265 22239 28187 22240
rect 21975 22112 22102 22128
rect 21975 21988 22079 22112
rect 21975 21972 22102 21988
rect 15946 21860 21868 21861
rect 15946 15940 15947 21860
rect 21867 15940 21868 21860
rect 15946 15939 21868 15940
rect 15656 15812 15783 15828
rect 15656 15688 15760 15812
rect 15656 15672 15783 15688
rect 9627 15560 15549 15561
rect 9627 9640 9628 15560
rect 15548 9640 15549 15560
rect 9627 9639 15549 9640
rect 9337 9512 9464 9528
rect 9337 9388 9441 9512
rect 9337 9372 9464 9388
rect 3308 9260 9230 9261
rect 3308 3340 3309 9260
rect 9229 3340 9230 9260
rect 3308 3339 9230 3340
rect 3018 3212 3145 3228
rect 3018 3088 3122 3212
rect 3018 3072 3145 3088
rect -3011 2960 2911 2961
rect -3011 -2960 -3010 2960
rect 2910 -2960 2911 2960
rect -3011 -2961 2911 -2960
rect -3301 -3088 -3174 -3072
rect -3301 -3212 -3197 -3088
rect -3301 -3228 -3174 -3212
rect -9330 -3340 -3408 -3339
rect -9330 -9260 -9329 -3340
rect -3409 -9260 -3408 -3340
rect -9330 -9261 -3408 -9260
rect -9620 -9388 -9493 -9372
rect -9620 -9512 -9516 -9388
rect -9620 -9528 -9493 -9512
rect -15649 -9640 -9727 -9639
rect -15649 -15560 -15648 -9640
rect -9728 -15560 -9727 -9640
rect -15649 -15561 -9727 -15560
rect -15939 -15688 -15812 -15672
rect -15939 -15812 -15835 -15688
rect -15939 -15828 -15812 -15812
rect -21968 -15940 -16046 -15939
rect -21968 -21860 -21967 -15940
rect -16047 -21860 -16046 -15940
rect -21968 -21861 -16046 -21860
rect -22258 -21988 -22131 -21972
rect -22258 -22112 -22154 -21988
rect -22258 -22128 -22131 -22112
rect -28287 -22240 -22365 -22239
rect -28287 -28160 -28286 -22240
rect -22366 -28160 -22365 -22240
rect -28287 -28161 -22365 -28160
rect -28577 -28288 -28450 -28272
rect -28577 -28412 -28473 -28288
rect -28577 -28428 -28450 -28412
rect -34606 -28540 -28684 -28539
rect -34606 -34460 -34605 -28540
rect -28685 -34460 -28684 -28540
rect -34606 -34461 -28684 -34460
rect -34896 -34588 -34769 -34572
rect -34896 -34712 -34792 -34588
rect -34896 -34728 -34769 -34712
rect -40925 -34840 -35003 -34839
rect -40925 -40760 -40924 -34840
rect -35004 -40760 -35003 -34840
rect -40925 -40761 -35003 -40760
rect -41215 -40888 -41088 -40872
rect -41215 -41012 -41111 -40888
rect -41215 -41028 -41088 -41012
rect -47244 -41140 -41322 -41139
rect -47244 -47060 -47243 -41140
rect -41323 -47060 -41322 -41140
rect -47244 -47061 -41322 -47060
rect -44335 -47250 -44231 -47061
rect -41215 -47172 -41168 -41028
rect -41104 -47172 -41088 -41028
rect -38016 -41139 -37912 -40761
rect -34896 -40872 -34849 -34728
rect -34785 -40872 -34769 -34728
rect -31697 -34839 -31593 -34461
rect -28577 -34572 -28530 -28428
rect -28466 -34572 -28450 -28428
rect -25378 -28539 -25274 -28161
rect -22258 -28272 -22211 -22128
rect -22147 -28272 -22131 -22128
rect -19059 -22239 -18955 -21861
rect -15939 -21972 -15892 -15828
rect -15828 -21972 -15812 -15828
rect -12740 -15939 -12636 -15561
rect -9620 -15672 -9573 -9528
rect -9509 -15672 -9493 -9528
rect -6421 -9639 -6317 -9261
rect -3301 -9372 -3254 -3228
rect -3190 -9372 -3174 -3228
rect -102 -3339 2 -2961
rect 3018 -3072 3065 3072
rect 3129 -3072 3145 3072
rect 6217 2961 6321 3339
rect 9337 3228 9384 9372
rect 9448 3228 9464 9372
rect 12536 9261 12640 9639
rect 15656 9528 15703 15672
rect 15767 9528 15783 15672
rect 18855 15561 18959 15939
rect 21975 15828 22022 21972
rect 22086 15828 22102 21972
rect 25174 21861 25278 22239
rect 28294 22128 28341 28272
rect 28405 22128 28421 28272
rect 31493 28161 31597 28539
rect 34613 28428 34660 34572
rect 34724 28428 34740 34572
rect 37812 34461 37916 34839
rect 40932 34728 40979 40872
rect 41043 34728 41059 40872
rect 44131 40761 44235 41139
rect 47251 41028 47298 47172
rect 47362 41028 47378 47172
rect 47251 41012 47378 41028
rect 47251 40888 47355 41012
rect 47251 40872 47378 40888
rect 41222 40760 47144 40761
rect 41222 34840 41223 40760
rect 47143 34840 47144 40760
rect 41222 34839 47144 34840
rect 40932 34712 41059 34728
rect 40932 34588 41036 34712
rect 40932 34572 41059 34588
rect 34903 34460 40825 34461
rect 34903 28540 34904 34460
rect 40824 28540 40825 34460
rect 34903 28539 40825 28540
rect 34613 28412 34740 28428
rect 34613 28288 34717 28412
rect 34613 28272 34740 28288
rect 28584 28160 34506 28161
rect 28584 22240 28585 28160
rect 34505 22240 34506 28160
rect 28584 22239 34506 22240
rect 28294 22112 28421 22128
rect 28294 21988 28398 22112
rect 28294 21972 28421 21988
rect 22265 21860 28187 21861
rect 22265 15940 22266 21860
rect 28186 15940 28187 21860
rect 22265 15939 28187 15940
rect 21975 15812 22102 15828
rect 21975 15688 22079 15812
rect 21975 15672 22102 15688
rect 15946 15560 21868 15561
rect 15946 9640 15947 15560
rect 21867 9640 21868 15560
rect 15946 9639 21868 9640
rect 15656 9512 15783 9528
rect 15656 9388 15760 9512
rect 15656 9372 15783 9388
rect 9627 9260 15549 9261
rect 9627 3340 9628 9260
rect 15548 3340 15549 9260
rect 9627 3339 15549 3340
rect 9337 3212 9464 3228
rect 9337 3088 9441 3212
rect 9337 3072 9464 3088
rect 3308 2960 9230 2961
rect 3308 -2960 3309 2960
rect 9229 -2960 9230 2960
rect 3308 -2961 9230 -2960
rect 3018 -3088 3145 -3072
rect 3018 -3212 3122 -3088
rect 3018 -3228 3145 -3212
rect -3011 -3340 2911 -3339
rect -3011 -9260 -3010 -3340
rect 2910 -9260 2911 -3340
rect -3011 -9261 2911 -9260
rect -3301 -9388 -3174 -9372
rect -3301 -9512 -3197 -9388
rect -3301 -9528 -3174 -9512
rect -9330 -9640 -3408 -9639
rect -9330 -15560 -9329 -9640
rect -3409 -15560 -3408 -9640
rect -9330 -15561 -3408 -15560
rect -9620 -15688 -9493 -15672
rect -9620 -15812 -9516 -15688
rect -9620 -15828 -9493 -15812
rect -15649 -15940 -9727 -15939
rect -15649 -21860 -15648 -15940
rect -9728 -21860 -9727 -15940
rect -15649 -21861 -9727 -21860
rect -15939 -21988 -15812 -21972
rect -15939 -22112 -15835 -21988
rect -15939 -22128 -15812 -22112
rect -21968 -22240 -16046 -22239
rect -21968 -28160 -21967 -22240
rect -16047 -28160 -16046 -22240
rect -21968 -28161 -16046 -28160
rect -22258 -28288 -22131 -28272
rect -22258 -28412 -22154 -28288
rect -22258 -28428 -22131 -28412
rect -28287 -28540 -22365 -28539
rect -28287 -34460 -28286 -28540
rect -22366 -34460 -22365 -28540
rect -28287 -34461 -22365 -34460
rect -28577 -34588 -28450 -34572
rect -28577 -34712 -28473 -34588
rect -28577 -34728 -28450 -34712
rect -34606 -34840 -28684 -34839
rect -34606 -40760 -34605 -34840
rect -28685 -40760 -28684 -34840
rect -34606 -40761 -28684 -40760
rect -34896 -40888 -34769 -40872
rect -34896 -41012 -34792 -40888
rect -34896 -41028 -34769 -41012
rect -40925 -41140 -35003 -41139
rect -40925 -47060 -40924 -41140
rect -35004 -47060 -35003 -41140
rect -40925 -47061 -35003 -47060
rect -41215 -47188 -41088 -47172
rect -41215 -47250 -41111 -47188
rect -38016 -47250 -37912 -47061
rect -34896 -47172 -34849 -41028
rect -34785 -47172 -34769 -41028
rect -31697 -41139 -31593 -40761
rect -28577 -40872 -28530 -34728
rect -28466 -40872 -28450 -34728
rect -25378 -34839 -25274 -34461
rect -22258 -34572 -22211 -28428
rect -22147 -34572 -22131 -28428
rect -19059 -28539 -18955 -28161
rect -15939 -28272 -15892 -22128
rect -15828 -28272 -15812 -22128
rect -12740 -22239 -12636 -21861
rect -9620 -21972 -9573 -15828
rect -9509 -21972 -9493 -15828
rect -6421 -15939 -6317 -15561
rect -3301 -15672 -3254 -9528
rect -3190 -15672 -3174 -9528
rect -102 -9639 2 -9261
rect 3018 -9372 3065 -3228
rect 3129 -9372 3145 -3228
rect 6217 -3339 6321 -2961
rect 9337 -3072 9384 3072
rect 9448 -3072 9464 3072
rect 12536 2961 12640 3339
rect 15656 3228 15703 9372
rect 15767 3228 15783 9372
rect 18855 9261 18959 9639
rect 21975 9528 22022 15672
rect 22086 9528 22102 15672
rect 25174 15561 25278 15939
rect 28294 15828 28341 21972
rect 28405 15828 28421 21972
rect 31493 21861 31597 22239
rect 34613 22128 34660 28272
rect 34724 22128 34740 28272
rect 37812 28161 37916 28539
rect 40932 28428 40979 34572
rect 41043 28428 41059 34572
rect 44131 34461 44235 34839
rect 47251 34728 47298 40872
rect 47362 34728 47378 40872
rect 47251 34712 47378 34728
rect 47251 34588 47355 34712
rect 47251 34572 47378 34588
rect 41222 34460 47144 34461
rect 41222 28540 41223 34460
rect 47143 28540 47144 34460
rect 41222 28539 47144 28540
rect 40932 28412 41059 28428
rect 40932 28288 41036 28412
rect 40932 28272 41059 28288
rect 34903 28160 40825 28161
rect 34903 22240 34904 28160
rect 40824 22240 40825 28160
rect 34903 22239 40825 22240
rect 34613 22112 34740 22128
rect 34613 21988 34717 22112
rect 34613 21972 34740 21988
rect 28584 21860 34506 21861
rect 28584 15940 28585 21860
rect 34505 15940 34506 21860
rect 28584 15939 34506 15940
rect 28294 15812 28421 15828
rect 28294 15688 28398 15812
rect 28294 15672 28421 15688
rect 22265 15560 28187 15561
rect 22265 9640 22266 15560
rect 28186 9640 28187 15560
rect 22265 9639 28187 9640
rect 21975 9512 22102 9528
rect 21975 9388 22079 9512
rect 21975 9372 22102 9388
rect 15946 9260 21868 9261
rect 15946 3340 15947 9260
rect 21867 3340 21868 9260
rect 15946 3339 21868 3340
rect 15656 3212 15783 3228
rect 15656 3088 15760 3212
rect 15656 3072 15783 3088
rect 9627 2960 15549 2961
rect 9627 -2960 9628 2960
rect 15548 -2960 15549 2960
rect 9627 -2961 15549 -2960
rect 9337 -3088 9464 -3072
rect 9337 -3212 9441 -3088
rect 9337 -3228 9464 -3212
rect 3308 -3340 9230 -3339
rect 3308 -9260 3309 -3340
rect 9229 -9260 9230 -3340
rect 3308 -9261 9230 -9260
rect 3018 -9388 3145 -9372
rect 3018 -9512 3122 -9388
rect 3018 -9528 3145 -9512
rect -3011 -9640 2911 -9639
rect -3011 -15560 -3010 -9640
rect 2910 -15560 2911 -9640
rect -3011 -15561 2911 -15560
rect -3301 -15688 -3174 -15672
rect -3301 -15812 -3197 -15688
rect -3301 -15828 -3174 -15812
rect -9330 -15940 -3408 -15939
rect -9330 -21860 -9329 -15940
rect -3409 -21860 -3408 -15940
rect -9330 -21861 -3408 -21860
rect -9620 -21988 -9493 -21972
rect -9620 -22112 -9516 -21988
rect -9620 -22128 -9493 -22112
rect -15649 -22240 -9727 -22239
rect -15649 -28160 -15648 -22240
rect -9728 -28160 -9727 -22240
rect -15649 -28161 -9727 -28160
rect -15939 -28288 -15812 -28272
rect -15939 -28412 -15835 -28288
rect -15939 -28428 -15812 -28412
rect -21968 -28540 -16046 -28539
rect -21968 -34460 -21967 -28540
rect -16047 -34460 -16046 -28540
rect -21968 -34461 -16046 -34460
rect -22258 -34588 -22131 -34572
rect -22258 -34712 -22154 -34588
rect -22258 -34728 -22131 -34712
rect -28287 -34840 -22365 -34839
rect -28287 -40760 -28286 -34840
rect -22366 -40760 -22365 -34840
rect -28287 -40761 -22365 -40760
rect -28577 -40888 -28450 -40872
rect -28577 -41012 -28473 -40888
rect -28577 -41028 -28450 -41012
rect -34606 -41140 -28684 -41139
rect -34606 -47060 -34605 -41140
rect -28685 -47060 -28684 -41140
rect -34606 -47061 -28684 -47060
rect -34896 -47188 -34769 -47172
rect -34896 -47250 -34792 -47188
rect -31697 -47250 -31593 -47061
rect -28577 -47172 -28530 -41028
rect -28466 -47172 -28450 -41028
rect -25378 -41139 -25274 -40761
rect -22258 -40872 -22211 -34728
rect -22147 -40872 -22131 -34728
rect -19059 -34839 -18955 -34461
rect -15939 -34572 -15892 -28428
rect -15828 -34572 -15812 -28428
rect -12740 -28539 -12636 -28161
rect -9620 -28272 -9573 -22128
rect -9509 -28272 -9493 -22128
rect -6421 -22239 -6317 -21861
rect -3301 -21972 -3254 -15828
rect -3190 -21972 -3174 -15828
rect -102 -15939 2 -15561
rect 3018 -15672 3065 -9528
rect 3129 -15672 3145 -9528
rect 6217 -9639 6321 -9261
rect 9337 -9372 9384 -3228
rect 9448 -9372 9464 -3228
rect 12536 -3339 12640 -2961
rect 15656 -3072 15703 3072
rect 15767 -3072 15783 3072
rect 18855 2961 18959 3339
rect 21975 3228 22022 9372
rect 22086 3228 22102 9372
rect 25174 9261 25278 9639
rect 28294 9528 28341 15672
rect 28405 9528 28421 15672
rect 31493 15561 31597 15939
rect 34613 15828 34660 21972
rect 34724 15828 34740 21972
rect 37812 21861 37916 22239
rect 40932 22128 40979 28272
rect 41043 22128 41059 28272
rect 44131 28161 44235 28539
rect 47251 28428 47298 34572
rect 47362 28428 47378 34572
rect 47251 28412 47378 28428
rect 47251 28288 47355 28412
rect 47251 28272 47378 28288
rect 41222 28160 47144 28161
rect 41222 22240 41223 28160
rect 47143 22240 47144 28160
rect 41222 22239 47144 22240
rect 40932 22112 41059 22128
rect 40932 21988 41036 22112
rect 40932 21972 41059 21988
rect 34903 21860 40825 21861
rect 34903 15940 34904 21860
rect 40824 15940 40825 21860
rect 34903 15939 40825 15940
rect 34613 15812 34740 15828
rect 34613 15688 34717 15812
rect 34613 15672 34740 15688
rect 28584 15560 34506 15561
rect 28584 9640 28585 15560
rect 34505 9640 34506 15560
rect 28584 9639 34506 9640
rect 28294 9512 28421 9528
rect 28294 9388 28398 9512
rect 28294 9372 28421 9388
rect 22265 9260 28187 9261
rect 22265 3340 22266 9260
rect 28186 3340 28187 9260
rect 22265 3339 28187 3340
rect 21975 3212 22102 3228
rect 21975 3088 22079 3212
rect 21975 3072 22102 3088
rect 15946 2960 21868 2961
rect 15946 -2960 15947 2960
rect 21867 -2960 21868 2960
rect 15946 -2961 21868 -2960
rect 15656 -3088 15783 -3072
rect 15656 -3212 15760 -3088
rect 15656 -3228 15783 -3212
rect 9627 -3340 15549 -3339
rect 9627 -9260 9628 -3340
rect 15548 -9260 15549 -3340
rect 9627 -9261 15549 -9260
rect 9337 -9388 9464 -9372
rect 9337 -9512 9441 -9388
rect 9337 -9528 9464 -9512
rect 3308 -9640 9230 -9639
rect 3308 -15560 3309 -9640
rect 9229 -15560 9230 -9640
rect 3308 -15561 9230 -15560
rect 3018 -15688 3145 -15672
rect 3018 -15812 3122 -15688
rect 3018 -15828 3145 -15812
rect -3011 -15940 2911 -15939
rect -3011 -21860 -3010 -15940
rect 2910 -21860 2911 -15940
rect -3011 -21861 2911 -21860
rect -3301 -21988 -3174 -21972
rect -3301 -22112 -3197 -21988
rect -3301 -22128 -3174 -22112
rect -9330 -22240 -3408 -22239
rect -9330 -28160 -9329 -22240
rect -3409 -28160 -3408 -22240
rect -9330 -28161 -3408 -28160
rect -9620 -28288 -9493 -28272
rect -9620 -28412 -9516 -28288
rect -9620 -28428 -9493 -28412
rect -15649 -28540 -9727 -28539
rect -15649 -34460 -15648 -28540
rect -9728 -34460 -9727 -28540
rect -15649 -34461 -9727 -34460
rect -15939 -34588 -15812 -34572
rect -15939 -34712 -15835 -34588
rect -15939 -34728 -15812 -34712
rect -21968 -34840 -16046 -34839
rect -21968 -40760 -21967 -34840
rect -16047 -40760 -16046 -34840
rect -21968 -40761 -16046 -40760
rect -22258 -40888 -22131 -40872
rect -22258 -41012 -22154 -40888
rect -22258 -41028 -22131 -41012
rect -28287 -41140 -22365 -41139
rect -28287 -47060 -28286 -41140
rect -22366 -47060 -22365 -41140
rect -28287 -47061 -22365 -47060
rect -28577 -47188 -28450 -47172
rect -28577 -47250 -28473 -47188
rect -25378 -47250 -25274 -47061
rect -22258 -47172 -22211 -41028
rect -22147 -47172 -22131 -41028
rect -19059 -41139 -18955 -40761
rect -15939 -40872 -15892 -34728
rect -15828 -40872 -15812 -34728
rect -12740 -34839 -12636 -34461
rect -9620 -34572 -9573 -28428
rect -9509 -34572 -9493 -28428
rect -6421 -28539 -6317 -28161
rect -3301 -28272 -3254 -22128
rect -3190 -28272 -3174 -22128
rect -102 -22239 2 -21861
rect 3018 -21972 3065 -15828
rect 3129 -21972 3145 -15828
rect 6217 -15939 6321 -15561
rect 9337 -15672 9384 -9528
rect 9448 -15672 9464 -9528
rect 12536 -9639 12640 -9261
rect 15656 -9372 15703 -3228
rect 15767 -9372 15783 -3228
rect 18855 -3339 18959 -2961
rect 21975 -3072 22022 3072
rect 22086 -3072 22102 3072
rect 25174 2961 25278 3339
rect 28294 3228 28341 9372
rect 28405 3228 28421 9372
rect 31493 9261 31597 9639
rect 34613 9528 34660 15672
rect 34724 9528 34740 15672
rect 37812 15561 37916 15939
rect 40932 15828 40979 21972
rect 41043 15828 41059 21972
rect 44131 21861 44235 22239
rect 47251 22128 47298 28272
rect 47362 22128 47378 28272
rect 47251 22112 47378 22128
rect 47251 21988 47355 22112
rect 47251 21972 47378 21988
rect 41222 21860 47144 21861
rect 41222 15940 41223 21860
rect 47143 15940 47144 21860
rect 41222 15939 47144 15940
rect 40932 15812 41059 15828
rect 40932 15688 41036 15812
rect 40932 15672 41059 15688
rect 34903 15560 40825 15561
rect 34903 9640 34904 15560
rect 40824 9640 40825 15560
rect 34903 9639 40825 9640
rect 34613 9512 34740 9528
rect 34613 9388 34717 9512
rect 34613 9372 34740 9388
rect 28584 9260 34506 9261
rect 28584 3340 28585 9260
rect 34505 3340 34506 9260
rect 28584 3339 34506 3340
rect 28294 3212 28421 3228
rect 28294 3088 28398 3212
rect 28294 3072 28421 3088
rect 22265 2960 28187 2961
rect 22265 -2960 22266 2960
rect 28186 -2960 28187 2960
rect 22265 -2961 28187 -2960
rect 21975 -3088 22102 -3072
rect 21975 -3212 22079 -3088
rect 21975 -3228 22102 -3212
rect 15946 -3340 21868 -3339
rect 15946 -9260 15947 -3340
rect 21867 -9260 21868 -3340
rect 15946 -9261 21868 -9260
rect 15656 -9388 15783 -9372
rect 15656 -9512 15760 -9388
rect 15656 -9528 15783 -9512
rect 9627 -9640 15549 -9639
rect 9627 -15560 9628 -9640
rect 15548 -15560 15549 -9640
rect 9627 -15561 15549 -15560
rect 9337 -15688 9464 -15672
rect 9337 -15812 9441 -15688
rect 9337 -15828 9464 -15812
rect 3308 -15940 9230 -15939
rect 3308 -21860 3309 -15940
rect 9229 -21860 9230 -15940
rect 3308 -21861 9230 -21860
rect 3018 -21988 3145 -21972
rect 3018 -22112 3122 -21988
rect 3018 -22128 3145 -22112
rect -3011 -22240 2911 -22239
rect -3011 -28160 -3010 -22240
rect 2910 -28160 2911 -22240
rect -3011 -28161 2911 -28160
rect -3301 -28288 -3174 -28272
rect -3301 -28412 -3197 -28288
rect -3301 -28428 -3174 -28412
rect -9330 -28540 -3408 -28539
rect -9330 -34460 -9329 -28540
rect -3409 -34460 -3408 -28540
rect -9330 -34461 -3408 -34460
rect -9620 -34588 -9493 -34572
rect -9620 -34712 -9516 -34588
rect -9620 -34728 -9493 -34712
rect -15649 -34840 -9727 -34839
rect -15649 -40760 -15648 -34840
rect -9728 -40760 -9727 -34840
rect -15649 -40761 -9727 -40760
rect -15939 -40888 -15812 -40872
rect -15939 -41012 -15835 -40888
rect -15939 -41028 -15812 -41012
rect -21968 -41140 -16046 -41139
rect -21968 -47060 -21967 -41140
rect -16047 -47060 -16046 -41140
rect -21968 -47061 -16046 -47060
rect -22258 -47188 -22131 -47172
rect -22258 -47250 -22154 -47188
rect -19059 -47250 -18955 -47061
rect -15939 -47172 -15892 -41028
rect -15828 -47172 -15812 -41028
rect -12740 -41139 -12636 -40761
rect -9620 -40872 -9573 -34728
rect -9509 -40872 -9493 -34728
rect -6421 -34839 -6317 -34461
rect -3301 -34572 -3254 -28428
rect -3190 -34572 -3174 -28428
rect -102 -28539 2 -28161
rect 3018 -28272 3065 -22128
rect 3129 -28272 3145 -22128
rect 6217 -22239 6321 -21861
rect 9337 -21972 9384 -15828
rect 9448 -21972 9464 -15828
rect 12536 -15939 12640 -15561
rect 15656 -15672 15703 -9528
rect 15767 -15672 15783 -9528
rect 18855 -9639 18959 -9261
rect 21975 -9372 22022 -3228
rect 22086 -9372 22102 -3228
rect 25174 -3339 25278 -2961
rect 28294 -3072 28341 3072
rect 28405 -3072 28421 3072
rect 31493 2961 31597 3339
rect 34613 3228 34660 9372
rect 34724 3228 34740 9372
rect 37812 9261 37916 9639
rect 40932 9528 40979 15672
rect 41043 9528 41059 15672
rect 44131 15561 44235 15939
rect 47251 15828 47298 21972
rect 47362 15828 47378 21972
rect 47251 15812 47378 15828
rect 47251 15688 47355 15812
rect 47251 15672 47378 15688
rect 41222 15560 47144 15561
rect 41222 9640 41223 15560
rect 47143 9640 47144 15560
rect 41222 9639 47144 9640
rect 40932 9512 41059 9528
rect 40932 9388 41036 9512
rect 40932 9372 41059 9388
rect 34903 9260 40825 9261
rect 34903 3340 34904 9260
rect 40824 3340 40825 9260
rect 34903 3339 40825 3340
rect 34613 3212 34740 3228
rect 34613 3088 34717 3212
rect 34613 3072 34740 3088
rect 28584 2960 34506 2961
rect 28584 -2960 28585 2960
rect 34505 -2960 34506 2960
rect 28584 -2961 34506 -2960
rect 28294 -3088 28421 -3072
rect 28294 -3212 28398 -3088
rect 28294 -3228 28421 -3212
rect 22265 -3340 28187 -3339
rect 22265 -9260 22266 -3340
rect 28186 -9260 28187 -3340
rect 22265 -9261 28187 -9260
rect 21975 -9388 22102 -9372
rect 21975 -9512 22079 -9388
rect 21975 -9528 22102 -9512
rect 15946 -9640 21868 -9639
rect 15946 -15560 15947 -9640
rect 21867 -15560 21868 -9640
rect 15946 -15561 21868 -15560
rect 15656 -15688 15783 -15672
rect 15656 -15812 15760 -15688
rect 15656 -15828 15783 -15812
rect 9627 -15940 15549 -15939
rect 9627 -21860 9628 -15940
rect 15548 -21860 15549 -15940
rect 9627 -21861 15549 -21860
rect 9337 -21988 9464 -21972
rect 9337 -22112 9441 -21988
rect 9337 -22128 9464 -22112
rect 3308 -22240 9230 -22239
rect 3308 -28160 3309 -22240
rect 9229 -28160 9230 -22240
rect 3308 -28161 9230 -28160
rect 3018 -28288 3145 -28272
rect 3018 -28412 3122 -28288
rect 3018 -28428 3145 -28412
rect -3011 -28540 2911 -28539
rect -3011 -34460 -3010 -28540
rect 2910 -34460 2911 -28540
rect -3011 -34461 2911 -34460
rect -3301 -34588 -3174 -34572
rect -3301 -34712 -3197 -34588
rect -3301 -34728 -3174 -34712
rect -9330 -34840 -3408 -34839
rect -9330 -40760 -9329 -34840
rect -3409 -40760 -3408 -34840
rect -9330 -40761 -3408 -40760
rect -9620 -40888 -9493 -40872
rect -9620 -41012 -9516 -40888
rect -9620 -41028 -9493 -41012
rect -15649 -41140 -9727 -41139
rect -15649 -47060 -15648 -41140
rect -9728 -47060 -9727 -41140
rect -15649 -47061 -9727 -47060
rect -15939 -47188 -15812 -47172
rect -15939 -47250 -15835 -47188
rect -12740 -47250 -12636 -47061
rect -9620 -47172 -9573 -41028
rect -9509 -47172 -9493 -41028
rect -6421 -41139 -6317 -40761
rect -3301 -40872 -3254 -34728
rect -3190 -40872 -3174 -34728
rect -102 -34839 2 -34461
rect 3018 -34572 3065 -28428
rect 3129 -34572 3145 -28428
rect 6217 -28539 6321 -28161
rect 9337 -28272 9384 -22128
rect 9448 -28272 9464 -22128
rect 12536 -22239 12640 -21861
rect 15656 -21972 15703 -15828
rect 15767 -21972 15783 -15828
rect 18855 -15939 18959 -15561
rect 21975 -15672 22022 -9528
rect 22086 -15672 22102 -9528
rect 25174 -9639 25278 -9261
rect 28294 -9372 28341 -3228
rect 28405 -9372 28421 -3228
rect 31493 -3339 31597 -2961
rect 34613 -3072 34660 3072
rect 34724 -3072 34740 3072
rect 37812 2961 37916 3339
rect 40932 3228 40979 9372
rect 41043 3228 41059 9372
rect 44131 9261 44235 9639
rect 47251 9528 47298 15672
rect 47362 9528 47378 15672
rect 47251 9512 47378 9528
rect 47251 9388 47355 9512
rect 47251 9372 47378 9388
rect 41222 9260 47144 9261
rect 41222 3340 41223 9260
rect 47143 3340 47144 9260
rect 41222 3339 47144 3340
rect 40932 3212 41059 3228
rect 40932 3088 41036 3212
rect 40932 3072 41059 3088
rect 34903 2960 40825 2961
rect 34903 -2960 34904 2960
rect 40824 -2960 40825 2960
rect 34903 -2961 40825 -2960
rect 34613 -3088 34740 -3072
rect 34613 -3212 34717 -3088
rect 34613 -3228 34740 -3212
rect 28584 -3340 34506 -3339
rect 28584 -9260 28585 -3340
rect 34505 -9260 34506 -3340
rect 28584 -9261 34506 -9260
rect 28294 -9388 28421 -9372
rect 28294 -9512 28398 -9388
rect 28294 -9528 28421 -9512
rect 22265 -9640 28187 -9639
rect 22265 -15560 22266 -9640
rect 28186 -15560 28187 -9640
rect 22265 -15561 28187 -15560
rect 21975 -15688 22102 -15672
rect 21975 -15812 22079 -15688
rect 21975 -15828 22102 -15812
rect 15946 -15940 21868 -15939
rect 15946 -21860 15947 -15940
rect 21867 -21860 21868 -15940
rect 15946 -21861 21868 -21860
rect 15656 -21988 15783 -21972
rect 15656 -22112 15760 -21988
rect 15656 -22128 15783 -22112
rect 9627 -22240 15549 -22239
rect 9627 -28160 9628 -22240
rect 15548 -28160 15549 -22240
rect 9627 -28161 15549 -28160
rect 9337 -28288 9464 -28272
rect 9337 -28412 9441 -28288
rect 9337 -28428 9464 -28412
rect 3308 -28540 9230 -28539
rect 3308 -34460 3309 -28540
rect 9229 -34460 9230 -28540
rect 3308 -34461 9230 -34460
rect 3018 -34588 3145 -34572
rect 3018 -34712 3122 -34588
rect 3018 -34728 3145 -34712
rect -3011 -34840 2911 -34839
rect -3011 -40760 -3010 -34840
rect 2910 -40760 2911 -34840
rect -3011 -40761 2911 -40760
rect -3301 -40888 -3174 -40872
rect -3301 -41012 -3197 -40888
rect -3301 -41028 -3174 -41012
rect -9330 -41140 -3408 -41139
rect -9330 -47060 -9329 -41140
rect -3409 -47060 -3408 -41140
rect -9330 -47061 -3408 -47060
rect -9620 -47188 -9493 -47172
rect -9620 -47250 -9516 -47188
rect -6421 -47250 -6317 -47061
rect -3301 -47172 -3254 -41028
rect -3190 -47172 -3174 -41028
rect -102 -41139 2 -40761
rect 3018 -40872 3065 -34728
rect 3129 -40872 3145 -34728
rect 6217 -34839 6321 -34461
rect 9337 -34572 9384 -28428
rect 9448 -34572 9464 -28428
rect 12536 -28539 12640 -28161
rect 15656 -28272 15703 -22128
rect 15767 -28272 15783 -22128
rect 18855 -22239 18959 -21861
rect 21975 -21972 22022 -15828
rect 22086 -21972 22102 -15828
rect 25174 -15939 25278 -15561
rect 28294 -15672 28341 -9528
rect 28405 -15672 28421 -9528
rect 31493 -9639 31597 -9261
rect 34613 -9372 34660 -3228
rect 34724 -9372 34740 -3228
rect 37812 -3339 37916 -2961
rect 40932 -3072 40979 3072
rect 41043 -3072 41059 3072
rect 44131 2961 44235 3339
rect 47251 3228 47298 9372
rect 47362 3228 47378 9372
rect 47251 3212 47378 3228
rect 47251 3088 47355 3212
rect 47251 3072 47378 3088
rect 41222 2960 47144 2961
rect 41222 -2960 41223 2960
rect 47143 -2960 47144 2960
rect 41222 -2961 47144 -2960
rect 40932 -3088 41059 -3072
rect 40932 -3212 41036 -3088
rect 40932 -3228 41059 -3212
rect 34903 -3340 40825 -3339
rect 34903 -9260 34904 -3340
rect 40824 -9260 40825 -3340
rect 34903 -9261 40825 -9260
rect 34613 -9388 34740 -9372
rect 34613 -9512 34717 -9388
rect 34613 -9528 34740 -9512
rect 28584 -9640 34506 -9639
rect 28584 -15560 28585 -9640
rect 34505 -15560 34506 -9640
rect 28584 -15561 34506 -15560
rect 28294 -15688 28421 -15672
rect 28294 -15812 28398 -15688
rect 28294 -15828 28421 -15812
rect 22265 -15940 28187 -15939
rect 22265 -21860 22266 -15940
rect 28186 -21860 28187 -15940
rect 22265 -21861 28187 -21860
rect 21975 -21988 22102 -21972
rect 21975 -22112 22079 -21988
rect 21975 -22128 22102 -22112
rect 15946 -22240 21868 -22239
rect 15946 -28160 15947 -22240
rect 21867 -28160 21868 -22240
rect 15946 -28161 21868 -28160
rect 15656 -28288 15783 -28272
rect 15656 -28412 15760 -28288
rect 15656 -28428 15783 -28412
rect 9627 -28540 15549 -28539
rect 9627 -34460 9628 -28540
rect 15548 -34460 15549 -28540
rect 9627 -34461 15549 -34460
rect 9337 -34588 9464 -34572
rect 9337 -34712 9441 -34588
rect 9337 -34728 9464 -34712
rect 3308 -34840 9230 -34839
rect 3308 -40760 3309 -34840
rect 9229 -40760 9230 -34840
rect 3308 -40761 9230 -40760
rect 3018 -40888 3145 -40872
rect 3018 -41012 3122 -40888
rect 3018 -41028 3145 -41012
rect -3011 -41140 2911 -41139
rect -3011 -47060 -3010 -41140
rect 2910 -47060 2911 -41140
rect -3011 -47061 2911 -47060
rect -3301 -47188 -3174 -47172
rect -3301 -47250 -3197 -47188
rect -102 -47250 2 -47061
rect 3018 -47172 3065 -41028
rect 3129 -47172 3145 -41028
rect 6217 -41139 6321 -40761
rect 9337 -40872 9384 -34728
rect 9448 -40872 9464 -34728
rect 12536 -34839 12640 -34461
rect 15656 -34572 15703 -28428
rect 15767 -34572 15783 -28428
rect 18855 -28539 18959 -28161
rect 21975 -28272 22022 -22128
rect 22086 -28272 22102 -22128
rect 25174 -22239 25278 -21861
rect 28294 -21972 28341 -15828
rect 28405 -21972 28421 -15828
rect 31493 -15939 31597 -15561
rect 34613 -15672 34660 -9528
rect 34724 -15672 34740 -9528
rect 37812 -9639 37916 -9261
rect 40932 -9372 40979 -3228
rect 41043 -9372 41059 -3228
rect 44131 -3339 44235 -2961
rect 47251 -3072 47298 3072
rect 47362 -3072 47378 3072
rect 47251 -3088 47378 -3072
rect 47251 -3212 47355 -3088
rect 47251 -3228 47378 -3212
rect 41222 -3340 47144 -3339
rect 41222 -9260 41223 -3340
rect 47143 -9260 47144 -3340
rect 41222 -9261 47144 -9260
rect 40932 -9388 41059 -9372
rect 40932 -9512 41036 -9388
rect 40932 -9528 41059 -9512
rect 34903 -9640 40825 -9639
rect 34903 -15560 34904 -9640
rect 40824 -15560 40825 -9640
rect 34903 -15561 40825 -15560
rect 34613 -15688 34740 -15672
rect 34613 -15812 34717 -15688
rect 34613 -15828 34740 -15812
rect 28584 -15940 34506 -15939
rect 28584 -21860 28585 -15940
rect 34505 -21860 34506 -15940
rect 28584 -21861 34506 -21860
rect 28294 -21988 28421 -21972
rect 28294 -22112 28398 -21988
rect 28294 -22128 28421 -22112
rect 22265 -22240 28187 -22239
rect 22265 -28160 22266 -22240
rect 28186 -28160 28187 -22240
rect 22265 -28161 28187 -28160
rect 21975 -28288 22102 -28272
rect 21975 -28412 22079 -28288
rect 21975 -28428 22102 -28412
rect 15946 -28540 21868 -28539
rect 15946 -34460 15947 -28540
rect 21867 -34460 21868 -28540
rect 15946 -34461 21868 -34460
rect 15656 -34588 15783 -34572
rect 15656 -34712 15760 -34588
rect 15656 -34728 15783 -34712
rect 9627 -34840 15549 -34839
rect 9627 -40760 9628 -34840
rect 15548 -40760 15549 -34840
rect 9627 -40761 15549 -40760
rect 9337 -40888 9464 -40872
rect 9337 -41012 9441 -40888
rect 9337 -41028 9464 -41012
rect 3308 -41140 9230 -41139
rect 3308 -47060 3309 -41140
rect 9229 -47060 9230 -41140
rect 3308 -47061 9230 -47060
rect 3018 -47188 3145 -47172
rect 3018 -47250 3122 -47188
rect 6217 -47250 6321 -47061
rect 9337 -47172 9384 -41028
rect 9448 -47172 9464 -41028
rect 12536 -41139 12640 -40761
rect 15656 -40872 15703 -34728
rect 15767 -40872 15783 -34728
rect 18855 -34839 18959 -34461
rect 21975 -34572 22022 -28428
rect 22086 -34572 22102 -28428
rect 25174 -28539 25278 -28161
rect 28294 -28272 28341 -22128
rect 28405 -28272 28421 -22128
rect 31493 -22239 31597 -21861
rect 34613 -21972 34660 -15828
rect 34724 -21972 34740 -15828
rect 37812 -15939 37916 -15561
rect 40932 -15672 40979 -9528
rect 41043 -15672 41059 -9528
rect 44131 -9639 44235 -9261
rect 47251 -9372 47298 -3228
rect 47362 -9372 47378 -3228
rect 47251 -9388 47378 -9372
rect 47251 -9512 47355 -9388
rect 47251 -9528 47378 -9512
rect 41222 -9640 47144 -9639
rect 41222 -15560 41223 -9640
rect 47143 -15560 47144 -9640
rect 41222 -15561 47144 -15560
rect 40932 -15688 41059 -15672
rect 40932 -15812 41036 -15688
rect 40932 -15828 41059 -15812
rect 34903 -15940 40825 -15939
rect 34903 -21860 34904 -15940
rect 40824 -21860 40825 -15940
rect 34903 -21861 40825 -21860
rect 34613 -21988 34740 -21972
rect 34613 -22112 34717 -21988
rect 34613 -22128 34740 -22112
rect 28584 -22240 34506 -22239
rect 28584 -28160 28585 -22240
rect 34505 -28160 34506 -22240
rect 28584 -28161 34506 -28160
rect 28294 -28288 28421 -28272
rect 28294 -28412 28398 -28288
rect 28294 -28428 28421 -28412
rect 22265 -28540 28187 -28539
rect 22265 -34460 22266 -28540
rect 28186 -34460 28187 -28540
rect 22265 -34461 28187 -34460
rect 21975 -34588 22102 -34572
rect 21975 -34712 22079 -34588
rect 21975 -34728 22102 -34712
rect 15946 -34840 21868 -34839
rect 15946 -40760 15947 -34840
rect 21867 -40760 21868 -34840
rect 15946 -40761 21868 -40760
rect 15656 -40888 15783 -40872
rect 15656 -41012 15760 -40888
rect 15656 -41028 15783 -41012
rect 9627 -41140 15549 -41139
rect 9627 -47060 9628 -41140
rect 15548 -47060 15549 -41140
rect 9627 -47061 15549 -47060
rect 9337 -47188 9464 -47172
rect 9337 -47250 9441 -47188
rect 12536 -47250 12640 -47061
rect 15656 -47172 15703 -41028
rect 15767 -47172 15783 -41028
rect 18855 -41139 18959 -40761
rect 21975 -40872 22022 -34728
rect 22086 -40872 22102 -34728
rect 25174 -34839 25278 -34461
rect 28294 -34572 28341 -28428
rect 28405 -34572 28421 -28428
rect 31493 -28539 31597 -28161
rect 34613 -28272 34660 -22128
rect 34724 -28272 34740 -22128
rect 37812 -22239 37916 -21861
rect 40932 -21972 40979 -15828
rect 41043 -21972 41059 -15828
rect 44131 -15939 44235 -15561
rect 47251 -15672 47298 -9528
rect 47362 -15672 47378 -9528
rect 47251 -15688 47378 -15672
rect 47251 -15812 47355 -15688
rect 47251 -15828 47378 -15812
rect 41222 -15940 47144 -15939
rect 41222 -21860 41223 -15940
rect 47143 -21860 47144 -15940
rect 41222 -21861 47144 -21860
rect 40932 -21988 41059 -21972
rect 40932 -22112 41036 -21988
rect 40932 -22128 41059 -22112
rect 34903 -22240 40825 -22239
rect 34903 -28160 34904 -22240
rect 40824 -28160 40825 -22240
rect 34903 -28161 40825 -28160
rect 34613 -28288 34740 -28272
rect 34613 -28412 34717 -28288
rect 34613 -28428 34740 -28412
rect 28584 -28540 34506 -28539
rect 28584 -34460 28585 -28540
rect 34505 -34460 34506 -28540
rect 28584 -34461 34506 -34460
rect 28294 -34588 28421 -34572
rect 28294 -34712 28398 -34588
rect 28294 -34728 28421 -34712
rect 22265 -34840 28187 -34839
rect 22265 -40760 22266 -34840
rect 28186 -40760 28187 -34840
rect 22265 -40761 28187 -40760
rect 21975 -40888 22102 -40872
rect 21975 -41012 22079 -40888
rect 21975 -41028 22102 -41012
rect 15946 -41140 21868 -41139
rect 15946 -47060 15947 -41140
rect 21867 -47060 21868 -41140
rect 15946 -47061 21868 -47060
rect 15656 -47188 15783 -47172
rect 15656 -47250 15760 -47188
rect 18855 -47250 18959 -47061
rect 21975 -47172 22022 -41028
rect 22086 -47172 22102 -41028
rect 25174 -41139 25278 -40761
rect 28294 -40872 28341 -34728
rect 28405 -40872 28421 -34728
rect 31493 -34839 31597 -34461
rect 34613 -34572 34660 -28428
rect 34724 -34572 34740 -28428
rect 37812 -28539 37916 -28161
rect 40932 -28272 40979 -22128
rect 41043 -28272 41059 -22128
rect 44131 -22239 44235 -21861
rect 47251 -21972 47298 -15828
rect 47362 -21972 47378 -15828
rect 47251 -21988 47378 -21972
rect 47251 -22112 47355 -21988
rect 47251 -22128 47378 -22112
rect 41222 -22240 47144 -22239
rect 41222 -28160 41223 -22240
rect 47143 -28160 47144 -22240
rect 41222 -28161 47144 -28160
rect 40932 -28288 41059 -28272
rect 40932 -28412 41036 -28288
rect 40932 -28428 41059 -28412
rect 34903 -28540 40825 -28539
rect 34903 -34460 34904 -28540
rect 40824 -34460 40825 -28540
rect 34903 -34461 40825 -34460
rect 34613 -34588 34740 -34572
rect 34613 -34712 34717 -34588
rect 34613 -34728 34740 -34712
rect 28584 -34840 34506 -34839
rect 28584 -40760 28585 -34840
rect 34505 -40760 34506 -34840
rect 28584 -40761 34506 -40760
rect 28294 -40888 28421 -40872
rect 28294 -41012 28398 -40888
rect 28294 -41028 28421 -41012
rect 22265 -41140 28187 -41139
rect 22265 -47060 22266 -41140
rect 28186 -47060 28187 -41140
rect 22265 -47061 28187 -47060
rect 21975 -47188 22102 -47172
rect 21975 -47250 22079 -47188
rect 25174 -47250 25278 -47061
rect 28294 -47172 28341 -41028
rect 28405 -47172 28421 -41028
rect 31493 -41139 31597 -40761
rect 34613 -40872 34660 -34728
rect 34724 -40872 34740 -34728
rect 37812 -34839 37916 -34461
rect 40932 -34572 40979 -28428
rect 41043 -34572 41059 -28428
rect 44131 -28539 44235 -28161
rect 47251 -28272 47298 -22128
rect 47362 -28272 47378 -22128
rect 47251 -28288 47378 -28272
rect 47251 -28412 47355 -28288
rect 47251 -28428 47378 -28412
rect 41222 -28540 47144 -28539
rect 41222 -34460 41223 -28540
rect 47143 -34460 47144 -28540
rect 41222 -34461 47144 -34460
rect 40932 -34588 41059 -34572
rect 40932 -34712 41036 -34588
rect 40932 -34728 41059 -34712
rect 34903 -34840 40825 -34839
rect 34903 -40760 34904 -34840
rect 40824 -40760 40825 -34840
rect 34903 -40761 40825 -40760
rect 34613 -40888 34740 -40872
rect 34613 -41012 34717 -40888
rect 34613 -41028 34740 -41012
rect 28584 -41140 34506 -41139
rect 28584 -47060 28585 -41140
rect 34505 -47060 34506 -41140
rect 28584 -47061 34506 -47060
rect 28294 -47188 28421 -47172
rect 28294 -47250 28398 -47188
rect 31493 -47250 31597 -47061
rect 34613 -47172 34660 -41028
rect 34724 -47172 34740 -41028
rect 37812 -41139 37916 -40761
rect 40932 -40872 40979 -34728
rect 41043 -40872 41059 -34728
rect 44131 -34839 44235 -34461
rect 47251 -34572 47298 -28428
rect 47362 -34572 47378 -28428
rect 47251 -34588 47378 -34572
rect 47251 -34712 47355 -34588
rect 47251 -34728 47378 -34712
rect 41222 -34840 47144 -34839
rect 41222 -40760 41223 -34840
rect 47143 -40760 47144 -34840
rect 41222 -40761 47144 -40760
rect 40932 -40888 41059 -40872
rect 40932 -41012 41036 -40888
rect 40932 -41028 41059 -41012
rect 34903 -41140 40825 -41139
rect 34903 -47060 34904 -41140
rect 40824 -47060 40825 -41140
rect 34903 -47061 40825 -47060
rect 34613 -47188 34740 -47172
rect 34613 -47250 34717 -47188
rect 37812 -47250 37916 -47061
rect 40932 -47172 40979 -41028
rect 41043 -47172 41059 -41028
rect 44131 -41139 44235 -40761
rect 47251 -40872 47298 -34728
rect 47362 -40872 47378 -34728
rect 47251 -40888 47378 -40872
rect 47251 -41012 47355 -40888
rect 47251 -41028 47378 -41012
rect 41222 -41140 47144 -41139
rect 41222 -47060 41223 -41140
rect 47143 -47060 47144 -41140
rect 41222 -47061 47144 -47060
rect 40932 -47188 41059 -47172
rect 40932 -47250 41036 -47188
rect 44131 -47250 44235 -47061
rect 47251 -47172 47298 -41028
rect 47362 -47172 47378 -41028
rect 47251 -47188 47378 -47172
rect 47251 -47250 47355 -47188
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX 41083 41000 47283 47200
string parameters w 30 l 30 val 1.822k carea 2.00 cperi 0.19 nx 15 ny 15 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
string library sky130
<< end >>
