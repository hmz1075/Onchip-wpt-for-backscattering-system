magic
tech sky130A
timestamp 1634546801
<< locali >>
rect 9136 11136 9269 11174
rect 9136 11053 9165 11136
rect 9228 11053 9269 11136
rect 9136 11024 9269 11053
rect 9245 10487 9334 10506
rect 9245 10434 9259 10487
rect 9304 10434 9334 10487
rect 9245 10423 9334 10434
<< viali >>
rect 9165 11053 9228 11136
rect 9259 10434 9304 10487
<< metal1 >>
rect 9136 11136 9269 11174
rect 9136 11053 9165 11136
rect 9228 11053 9269 11136
rect 9136 11024 9269 11053
rect 10232 10616 10419 11078
rect 12908 10558 13160 11114
rect 15371 10591 15553 11111
rect 9245 10487 9334 10506
rect 9245 10434 9259 10487
rect 9304 10434 9334 10487
rect 9245 10423 9334 10434
<< via1 >>
rect 9259 10434 9304 10487
<< metal2 >>
rect 8638 19074 9280 19189
rect 18393 11218 19133 11221
rect 18331 11201 19133 11218
rect 18331 11110 18910 11201
rect 19111 11110 19133 11201
rect 18331 11089 19133 11110
rect 9245 10487 9334 10506
rect 9245 10434 9259 10487
rect 9304 10434 9334 10487
rect 9245 10423 9334 10434
rect 18331 10415 18585 11089
rect 8621 2131 20244 2175
rect 8621 2007 19781 2131
rect 20161 2007 20244 2131
rect 8621 1972 20244 2007
<< via2 >>
rect 18910 11110 19111 11201
rect 19781 2007 20161 2131
<< metal3 >>
rect 18890 11201 19136 11221
rect 18890 11110 18910 11201
rect 19111 11110 19136 11201
rect 18890 11086 19136 11110
<< via3 >>
rect 18910 11110 19111 11201
<< metal4 >>
rect 19675 11243 21189 11483
rect 18890 11201 21189 11243
rect 18890 11110 18910 11201
rect 19111 11110 21189 11201
rect 18890 11078 21189 11110
rect 19645 10828 21189 11078
use recitifer_layout  recitifer_layout_0
timestamp 1634373541
transform 1 0 465 0 1 14659
box -455 -14659 8736 4737
use cap225_layout  cap225_layout_0
timestamp 1634294201
transform 1 0 64697 0 1 44933
box -45016 -44796 3719 4460
use pmos40  pmos40_0
timestamp 1634376359
transform 1 0 9140 0 -1 19362
box 0 0 9454 8332
use pmos40  pmos40_1
timestamp 1634376359
transform 1 0 9203 0 -1 10682
box 0 0 9454 8332
<< labels >>
rlabel metal4 19242 11193 19242 11193 1 VIN2
rlabel metal2 9030 19129 9030 19129 1 VIN1
rlabel metal2 19358 2062 19358 2062 1 VSS
rlabel metal1 13066 10807 13066 10807 1 VOUT_C
rlabel space 9236 2465 9236 2465 1 VOUT
<< end >>
