**.subckt PICOOAYOUT
XM1 VINP VINN GND GND sky130_fd_pr__nfet_01v8_lvt L=0.35 W=80 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=20 m=20 
XM2 VINN VINP GND GND sky130_fd_pr__nfet_01v8_lvt L=0.35 W=80 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=20 m=20 
XM4 VIN1 VINP VINN VINN sky130_fd_pr__pfet_01v8_lvt L=0.35 W=80 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=20 m=20 
XM3 VIN1 VINN VINP VINP sky130_fd_pr__pfet_01v8_lvt L=0.35 W=80 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=20 m=20 
VSIN2 VINP VINN SIN(0 0.5 200MEG 0 0)
XM5 VOUT VOUT_C VIN1 VOUT sky130_fd_pr__pfet_01v8_lvt L=0.35 W=80 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=40 m=40 
XM6 VIN1 net2 net3 VIN1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=50 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM7 net4 VOUT net2 VSS sky130_fd_pr__nfet_01v8_lvt L=0.350 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM8 net4 VIN1 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.35 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM9 net2 net3 VIN1 VIN1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=50 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM10 VOUT_C net2 VOUT VIN1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=50 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM11 VOUT_C VOUT net5 VSS sky130_fd_pr__nfet_01v8_lvt L=0.35 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM12 net3 VIN1 net4 VSS sky130_fd_pr__nfet_01v8_lvt L=0.35 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM13 net5 VIN1 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.35 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
V1 VSS GND 0
VSIN1 __UNCONNECTED_PIN__0 GND 0
VSIN3 net1 GND 0
XM14 VREC VOUT_C VOUT VOUT sky130_fd_pr__pfet_01v8_lvt L=0.35 W=80 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=40 m=40 
XC3 VOUT net1 sky130_fd_pr__cap_mim_m3_1 W=30 L=30 MF=225 m=225
**** begin user architecture code


	.control
	save all
	tran 1ns 20us
	Let PIN1= AVG(VINP*(i(VSIN2)))
	Let PIN2= AVG(VINN*(i(VSIN2)))
	Let PIN=PIN2+PIN2
	Let POUT1= AVG(VOUT*(i(VSIN3)))
	Let POUT2= AVG(VOUT*(i(VSIN1)))
	Let POUT=POUT1+POUT2

	Let EFF=(POUT/PIN)

	*plot VOUT VIN1
	*plot PIN
	plot POUT
	plot VOUT
	*plot POUT1
	*plot POUT2
	plot EFF
	*plot VOUT_C
	plot VREC



	*plot POUT


.endc


 ** manual skywater pdks install (with patches applied)
* .lib /home/shahid/open_pdks/sky130A/libs.tech/ngspice/models/sky130.lib.spice tt

** opencircuitdesign pdks install
.lib /home/shahid/open_pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt

.param mc_mm_switch=0
.param mc_pr_switch=0

**** end user architecture code
**.ends
.GLOBAL GND
** flattened .save nodes
.end
