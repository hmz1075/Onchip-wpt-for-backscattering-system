magic
tech sky130A
magscale 1 2
timestamp 1634724870
<< metal3 >>
rect -48352 6826 -39104 7354
rect -87990 6736 -39104 6826
rect -87990 -41534 8182 6736
rect -87990 -83286 -44124 -41534
rect -43036 -42600 8182 -41534
<< metal4 >>
rect -85248 7686 5658 10526
rect -43640 7016 -40250 7686
rect -43640 5666 -38556 7016
rect -35080 6600 4654 7686
rect -35080 6220 4762 6600
rect -85910 2668 -38556 5666
rect -38794 1668 -38556 2668
rect -43640 -46 -38556 1668
rect -86194 -3044 -38556 -46
rect -43640 -5972 -38556 -3044
rect -86194 -8970 -38556 -5972
rect -43640 -12326 -38556 -8970
rect -86480 -15324 -38556 -12326
rect -43640 -18464 -38556 -15324
rect -86410 -21462 -38556 -18464
rect -43640 -24318 -38556 -21462
rect -86266 -27316 -38556 -24318
rect -43640 -29886 -38556 -27316
rect -87122 -32884 -38556 -29886
rect -43640 -36526 -38556 -32884
rect -86338 -39524 -38556 -36526
rect -43640 -42666 -38556 -39524
rect -86480 -43664 -38556 -42666
rect -34968 -43664 -32492 6220
rect -28078 -43664 -25602 6220
rect -22390 -43664 -19914 6220
rect -16140 -43664 -13664 6220
rect -10292 -43664 -7816 6220
rect -4202 -43664 -1726 6220
rect 1886 -43664 4762 6220
rect -86480 -45664 5972 -43664
rect -43640 -46446 5972 -45664
rect -43640 -48806 -40250 -46446
rect -86766 -51804 -39650 -48806
rect -43640 -54374 -40250 -51804
rect -87122 -57372 -40006 -54374
rect -43640 -60656 -40250 -57372
rect -86980 -63654 -39864 -60656
rect -43640 -66154 -40250 -63654
rect -86908 -69152 -39792 -66154
rect -43640 -72078 -40250 -69152
rect -86766 -75076 -39650 -72078
rect -43640 -78432 -40250 -75076
rect -87266 -81430 -40150 -78432
rect -43640 -83672 -40250 -81430
use sky130_fd_pr__cap_mim_m3_1_V8VXPF  sky130_fd_pr__cap_mim_m3_1_V8VXPF_0
timestamp 1634724870
transform 0 1 -66286 -1 0 -38028
box -45133 -21000 45132 21000
use sky130_fd_pr__cap_mim_m3_1_NBPZFR  sky130_fd_pr__cap_mim_m3_1_NBPZFR_0
timestamp 1634546801
transform 1 0 -18247 0 1 -18230
box -24306 -24240 24306 24240
<< labels >>
rlabel metal3 -37108 6230 -37108 6230 1 VOUT
rlabel metal4 -38992 -44062 -38992 -44062 1 VIN
<< end >>
