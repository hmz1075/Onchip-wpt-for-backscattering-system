magic
tech sky130A
timestamp 1634734342
<< metal2 >>
rect 24917 3040 138308 3074
rect 24917 2453 200724 3040
rect 137028 2417 200724 2453
<< metal3 >>
rect -89205 161220 -82473 162258
rect -89205 156191 -87923 161220
rect -83540 156191 -82473 161220
rect -89205 46976 -82473 156191
rect -89192 46679 -82482 46976
rect 137095 46796 199770 47099
rect -89502 46628 -57922 46679
rect -89502 43587 2738 46628
rect 74514 43845 199770 46796
rect 74514 43797 137695 43845
rect -89502 43362 -57922 43587
<< via3 >>
rect -87923 156191 -83540 161220
<< metal4 >>
rect -89367 161220 -82595 162415
rect -89367 156191 -87923 161220
rect -83540 156191 -82595 161220
rect -89367 155095 -82595 156191
rect 790 50827 1333 54376
rect 2744 50827 4464 54376
rect 790 50777 4464 50827
rect 939 46511 3097 50777
rect 137433 25968 200196 26080
rect 137433 25909 200979 25968
rect 72834 23348 200979 25909
rect 137433 23296 200979 23348
<< via4 >>
rect -87923 156191 -83540 161220
rect 1333 50827 2744 54376
<< metal5 >>
rect -89367 161220 -82595 162415
rect -89367 156191 -87923 161220
rect -83540 156191 -82595 161220
rect -89367 155095 -82595 156191
rect -64449 56500 -58954 56907
rect -64449 54376 7599 56500
rect -64449 51005 1333 54376
rect -64449 -13717 -58954 51005
rect 66 50827 1333 51005
rect 2744 51005 7599 54376
rect 2744 50827 4799 51005
rect 66 50620 4799 50827
rect 66 50534 3648 50620
use INDUCTOR_layout  INDUCTOR_layout_0
timestamp 1634733432
transform 1 0 -483261 0 -1 1593239
box 394000 1431000 683000 1631000
use FINAL_without_ind  FINAL_without_ind_0
timestamp 1634725508
transform 1 0 6485 0 1 0
box -28962 0 68406 49393
<< labels >>
rlabel metal2 137761 2661 137761 2705 1 VOUT
rlabel metal3 137213 45270 137213 45270 1 VSS
rlabel metal4 137582 24671 137582 24671 1 VOUT_RECT
flabel metal3 137369 45269 137369 45269 0 FreeSans 80000 0 0 0 VSS
flabel metal4 138081 24967 138081 24967 0 FreeSans 80000 0 0 0 VOUT_RECT
flabel metal2 137725 2884 137725 2884 0 FreeSans 80000 0 0 0 VOUT
<< end >>
