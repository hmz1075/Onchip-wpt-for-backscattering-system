magic
tech sky130A
magscale 1 2
timestamp 1634288453
<< locali >>
rect -44 8214 9194 8270
rect -44 8212 5634 8214
rect -44 8210 3784 8212
rect -44 8208 1014 8210
rect -44 8198 90 8208
rect 232 8206 1014 8208
rect 232 8198 548 8206
rect 690 8198 1014 8206
rect 1156 8204 1936 8210
rect 1156 8198 1476 8204
rect 1618 8198 1936 8204
rect 2078 8208 2862 8210
rect 2078 8198 2398 8208
rect 2540 8198 2862 8208
rect 3004 8198 3324 8210
rect 3466 8198 3784 8210
rect 3926 8210 5634 8212
rect 3926 8206 4708 8210
rect 3926 8198 4246 8206
rect 4388 8198 4708 8206
rect 4850 8198 5168 8210
rect 5310 8198 5634 8210
rect 5776 8198 6096 8214
rect 6238 8212 9194 8214
rect 6238 8198 6556 8212
rect 6698 8210 7942 8212
rect 6698 8208 7482 8210
rect 6698 8198 7018 8208
rect 7160 8198 7482 8208
rect 7624 8198 7942 8210
rect 8084 8198 8404 8212
rect 8546 8198 8868 8212
rect 9010 8198 9194 8212
rect -52 -8038 88 -8028
rect 230 -8036 550 -8028
rect 692 -8036 1014 -8028
rect 1156 -8034 1478 -8028
rect 1620 -8034 1936 -8028
rect 2078 -8034 2400 -8028
rect 1156 -8036 2400 -8034
rect 2542 -8032 2862 -8028
rect 3004 -8032 3322 -8028
rect 2542 -8034 3322 -8032
rect 3464 -8034 3786 -8028
rect 3928 -8034 4250 -8028
rect 2542 -8036 4250 -8034
rect 4392 -8034 4712 -8028
rect 4854 -8034 5172 -8028
rect 5314 -8034 5636 -8028
rect 5778 -8032 6096 -8028
rect 6238 -8032 6558 -8028
rect 5778 -8034 6558 -8032
rect 4392 -8036 6558 -8034
rect 6700 -8032 7022 -8028
rect 7164 -8032 7484 -8028
rect 7626 -8032 7942 -8028
rect 6700 -8034 7942 -8032
rect 8084 -8034 8402 -8028
rect 8544 -8034 8868 -8028
rect 9010 -8034 9158 -8028
rect 6700 -8036 9158 -8034
rect 230 -8038 9158 -8036
rect -52 -8116 9158 -8038
<< metal1 >>
rect 120 8118 9114 8286
rect -166 8050 112 8072
rect -166 7982 -130 8050
rect 20 7982 112 8050
rect -166 7954 112 7982
rect 430 8050 572 8072
rect 430 7972 446 8050
rect 526 7972 572 8050
rect 430 7954 572 7972
rect 890 7990 926 8068
rect 1006 7990 1034 8068
rect 890 7952 1034 7990
rect 1354 8060 1496 8074
rect 1354 7982 1374 8060
rect 1454 7982 1496 8060
rect 1354 7950 1496 7982
rect 1806 8052 1962 8074
rect 1806 7974 1822 8052
rect 1902 7974 1962 8052
rect 1806 7940 1962 7974
rect 2278 8062 2422 8074
rect 2278 7984 2290 8062
rect 2370 7984 2422 8062
rect 2278 7942 2422 7984
rect 2732 8062 2884 8078
rect 2732 7984 2750 8062
rect 2830 7984 2884 8062
rect 2732 7940 2884 7984
rect 3200 8058 3350 8080
rect 3200 7980 3218 8058
rect 3298 7980 3350 8058
rect 3200 7942 3350 7980
rect 3702 8038 3808 8084
rect 3702 7960 3720 8038
rect 3800 7960 3808 8038
rect 3702 7942 3808 7960
rect 4122 8054 4272 8084
rect 4122 7976 4150 8054
rect 4230 7976 4272 8054
rect 4122 7950 4272 7976
rect 4582 8062 4732 8078
rect 4582 7984 4602 8062
rect 4682 7984 4732 8062
rect 4582 7954 4732 7984
rect 5082 8048 5196 8084
rect 5162 7970 5196 8048
rect 5082 7950 5196 7970
rect 5512 8046 5654 8086
rect 5512 7968 5528 8046
rect 5608 7968 5654 8046
rect 5970 8068 6118 8084
rect 5970 7990 6010 8068
rect 6090 7990 6118 8068
rect 5970 7968 6118 7990
rect 6434 8062 6574 8086
rect 6434 7984 6454 8062
rect 6534 7984 6574 8062
rect 5512 7948 5654 7968
rect 6434 7966 6574 7984
rect 6896 8062 7040 8082
rect 6896 7984 6912 8062
rect 6992 7984 7040 8062
rect 6896 7962 7040 7984
rect 7392 8056 7504 8070
rect 7392 7978 7404 8056
rect 7484 7978 7504 8056
rect 7392 7962 7504 7978
rect 7854 8064 7964 8066
rect 7854 7986 7864 8064
rect 7944 7986 7964 8064
rect 7854 7966 7964 7986
rect 8316 7996 8328 8074
rect 8408 7996 8426 8074
rect 8316 7964 8426 7996
rect 8750 8062 8888 8072
rect 8750 7984 8754 8062
rect 8834 7984 8888 8062
rect 8750 7964 8888 7984
rect 204 -7818 316 -7790
rect 204 -7896 230 -7818
rect 310 -7896 316 -7818
rect 204 -7906 316 -7896
rect 666 -7804 788 -7788
rect 666 -7882 692 -7804
rect 772 -7882 788 -7804
rect 666 -7906 788 -7882
rect 1118 -7804 1242 -7786
rect 1118 -7882 1148 -7804
rect 1228 -7882 1242 -7804
rect 1118 -7916 1242 -7882
rect 1590 -7808 1708 -7780
rect 1590 -7886 1612 -7808
rect 1692 -7886 1708 -7808
rect 1590 -7916 1708 -7886
rect 2046 -7800 2166 -7782
rect 2046 -7878 2068 -7800
rect 2148 -7878 2166 -7800
rect 2046 -7916 2166 -7878
rect 2504 -7810 2632 -7776
rect 2504 -7888 2536 -7810
rect 2616 -7888 2632 -7810
rect 2504 -7916 2632 -7888
rect 2964 -7790 3092 -7770
rect 2964 -7868 3010 -7790
rect 3090 -7868 3092 -7790
rect 2964 -7918 3092 -7868
rect 3430 -7802 3558 -7774
rect 3430 -7880 3460 -7802
rect 3540 -7880 3558 -7802
rect 3430 -7918 3558 -7880
rect 3894 -7800 4018 -7770
rect 3894 -7878 3932 -7800
rect 4012 -7878 4018 -7800
rect 3894 -7920 4018 -7878
rect 4354 -7792 4484 -7768
rect 4354 -7870 4396 -7792
rect 4476 -7870 4484 -7792
rect 4354 -7916 4484 -7870
rect 4814 -7792 4942 -7760
rect 4814 -7870 4858 -7792
rect 4938 -7870 4942 -7792
rect 4814 -7918 4942 -7870
rect 5292 -7782 5434 -7766
rect 5292 -7860 5310 -7782
rect 5390 -7860 5434 -7782
rect 5292 -7902 5434 -7860
rect 5752 -7798 5898 -7764
rect 5752 -7876 5768 -7798
rect 5848 -7876 5898 -7798
rect 5752 -7920 5898 -7876
rect 6214 -7786 6362 -7768
rect 6214 -7864 6240 -7786
rect 6320 -7864 6362 -7786
rect 6214 -7902 6362 -7864
rect 6674 -7780 6824 -7764
rect 6674 -7858 6734 -7780
rect 6814 -7858 6824 -7780
rect 6674 -7906 6824 -7858
rect 7136 -7774 7290 -7766
rect 7136 -7852 7180 -7774
rect 7260 -7852 7290 -7774
rect 7136 -7920 7290 -7852
rect 7600 -7780 7744 -7772
rect 7600 -7858 7644 -7780
rect 7724 -7858 7744 -7780
rect 7600 -7902 7744 -7858
rect 8060 -7782 8216 -7768
rect 8060 -7860 8106 -7782
rect 8186 -7860 8216 -7782
rect 8060 -7900 8216 -7860
rect 8520 -7784 8670 -7778
rect 8520 -7862 8564 -7784
rect 8644 -7862 8670 -7784
rect 8520 -7902 8670 -7862
rect 8986 -7788 9138 -7762
rect 8986 -7866 9024 -7788
rect 9104 -7866 9138 -7788
rect 8986 -7906 9138 -7866
rect 114 -8222 9138 -7950
<< via1 >>
rect -130 7982 20 8050
rect 446 7972 526 8050
rect 926 7990 1006 8068
rect 1374 7982 1454 8060
rect 1822 7974 1902 8052
rect 2290 7984 2370 8062
rect 2750 7984 2830 8062
rect 3218 7980 3298 8058
rect 3720 7960 3800 8038
rect 4150 7976 4230 8054
rect 4602 7984 4682 8062
rect 5082 7970 5162 8048
rect 5528 7968 5608 8046
rect 6010 7990 6090 8068
rect 6454 7984 6534 8062
rect 6912 7984 6992 8062
rect 7404 7978 7484 8056
rect 7864 7986 7944 8064
rect 8328 7996 8408 8074
rect 8754 7984 8834 8062
rect 230 -7896 310 -7818
rect 692 -7882 772 -7804
rect 1148 -7882 1228 -7804
rect 1612 -7886 1692 -7808
rect 2068 -7878 2148 -7800
rect 2536 -7888 2616 -7810
rect 3010 -7868 3090 -7790
rect 3460 -7880 3540 -7802
rect 3932 -7878 4012 -7800
rect 4396 -7870 4476 -7792
rect 4858 -7870 4938 -7792
rect 5310 -7860 5390 -7782
rect 5768 -7876 5848 -7798
rect 6240 -7864 6320 -7786
rect 6734 -7858 6814 -7780
rect 7180 -7852 7260 -7774
rect 7644 -7858 7724 -7780
rect 8106 -7860 8186 -7782
rect 8564 -7862 8644 -7784
rect 9024 -7866 9104 -7788
<< metal2 >>
rect 2278 8084 2884 8088
rect 4602 8086 5194 8088
rect 6026 8086 6576 8088
rect 3200 8084 3810 8086
rect 2278 8080 4274 8084
rect 4602 8080 7040 8086
rect -166 8072 572 8078
rect 2278 8074 7040 8080
rect 1398 8072 7040 8074
rect 7864 8082 8426 8086
rect 7864 8074 8890 8082
rect 7864 8072 8328 8074
rect -166 8068 8328 8072
rect -166 8050 926 8068
rect -166 7982 -130 8050
rect 20 7982 446 8050
rect -166 7972 446 7982
rect 526 7990 926 8050
rect 1006 8062 6010 8068
rect 1006 8060 2290 8062
rect 1006 7990 1374 8060
rect 526 7982 1374 7990
rect 1454 8052 2290 8060
rect 1454 7982 1822 8052
rect 526 7974 1822 7982
rect 1902 7984 2290 8052
rect 2370 7984 2750 8062
rect 2830 8058 4602 8062
rect 2830 7984 3218 8058
rect 1902 7980 3218 7984
rect 3298 8054 4602 8058
rect 3298 8038 4150 8054
rect 3298 7980 3720 8038
rect 1902 7974 3720 7980
rect 526 7972 3720 7974
rect -166 7960 3720 7972
rect 3800 7976 4150 8038
rect 4230 7984 4602 8054
rect 4682 8048 6010 8062
rect 4682 7984 5082 8048
rect 4230 7976 5082 7984
rect 3800 7970 5082 7976
rect 5162 8046 6010 8048
rect 5162 7970 5528 8046
rect 3800 7968 5528 7970
rect 5608 7990 6010 8046
rect 6090 8064 8328 8068
rect 6090 8062 7864 8064
rect 6090 7990 6454 8062
rect 5608 7984 6454 7990
rect 6534 7984 6912 8062
rect 6992 8056 7864 8062
rect 6992 7984 7404 8056
rect 5608 7978 7404 7984
rect 7484 7986 7864 8056
rect 7944 7996 8328 8064
rect 8408 8062 8890 8074
rect 8408 7996 8754 8062
rect 7944 7986 8754 7996
rect 7484 7984 8754 7986
rect 8834 7984 8890 8062
rect 7484 7978 8890 7984
rect 5608 7968 8890 7978
rect 3800 7960 5656 7968
rect 6026 7964 8890 7968
rect 6432 7962 8426 7964
rect 6432 7960 7506 7962
rect -166 7954 5656 7960
rect 928 7952 5656 7954
rect 928 7950 4274 7952
rect 1398 7948 4274 7950
rect 5084 7948 5656 7952
rect 1398 7942 3810 7948
rect 1910 7940 2884 7942
rect 2278 7938 2884 7940
rect 3200 7938 3810 7942
rect 6212 -7762 6826 -7760
rect 4360 -7766 7290 -7762
rect 8522 -7764 9136 -7760
rect 8064 -7766 9136 -7764
rect 3892 -7768 9136 -7766
rect 3428 -7770 9136 -7768
rect 2962 -7774 9136 -7770
rect 2502 -7778 7180 -7774
rect 1588 -7780 7180 -7778
rect 1588 -7782 6734 -7780
rect 1126 -7786 5310 -7782
rect 692 -7790 5310 -7786
rect -308 -7800 3010 -7790
rect -308 -7804 2068 -7800
rect -308 -7818 692 -7804
rect -308 -7896 230 -7818
rect 310 -7882 692 -7818
rect 772 -7882 1148 -7804
rect 1228 -7808 2068 -7804
rect 1228 -7882 1612 -7808
rect 310 -7886 1612 -7882
rect 1692 -7878 2068 -7808
rect 2148 -7810 3010 -7800
rect 2148 -7878 2536 -7810
rect 1692 -7886 2536 -7878
rect 310 -7888 2536 -7886
rect 2616 -7868 3010 -7810
rect 3090 -7792 5310 -7790
rect 3090 -7800 4396 -7792
rect 3090 -7802 3932 -7800
rect 3090 -7868 3460 -7802
rect 2616 -7880 3460 -7868
rect 3540 -7878 3932 -7802
rect 4012 -7870 4396 -7800
rect 4476 -7870 4858 -7792
rect 4938 -7860 5310 -7792
rect 5390 -7786 6734 -7782
rect 5390 -7798 6240 -7786
rect 5390 -7860 5768 -7798
rect 4938 -7870 5768 -7860
rect 4012 -7876 5768 -7870
rect 5848 -7864 6240 -7798
rect 6320 -7858 6734 -7786
rect 6814 -7852 7180 -7780
rect 7260 -7780 9136 -7774
rect 7260 -7852 7644 -7780
rect 6814 -7858 7644 -7852
rect 7724 -7782 9136 -7780
rect 7724 -7858 8106 -7782
rect 6320 -7860 8106 -7858
rect 8186 -7784 9136 -7782
rect 8186 -7860 8564 -7784
rect 6320 -7862 8564 -7860
rect 8644 -7788 9136 -7784
rect 8644 -7862 9024 -7788
rect 6320 -7864 9024 -7862
rect 5848 -7866 9024 -7864
rect 9104 -7866 9136 -7788
rect 5848 -7876 9136 -7866
rect 4012 -7878 9136 -7876
rect 3540 -7880 9136 -7878
rect 2616 -7888 9136 -7880
rect 310 -7896 9136 -7888
rect -308 -7906 9136 -7896
rect 692 -7916 9136 -7906
rect 2036 -7918 9136 -7916
rect 2502 -7920 9136 -7918
rect 3428 -7924 4018 -7920
rect 4360 -7922 9136 -7920
rect 4814 -7924 5900 -7922
rect 7132 -7924 9136 -7922
rect 4814 -7926 5438 -7924
use sky130_fd_pr__nfet_01v8_lvt_BPY4AF  sky130_fd_pr__nfet_01v8_lvt_BPY4AF_0
array 19 0 462 0 0 16420
timestamp 1634288381
transform 1 0 159 0 1 85
box -231 -8210 231 8210
<< labels >>
rlabel locali -14 8224 -14 8224 1 B
rlabel metal1 242 8152 242 8152 1 G
rlabel metal2 -142 8020 -142 8020 1 D
rlabel metal2 -204 -7864 -204 -7864 1 S
<< end >>
